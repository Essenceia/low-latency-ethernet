//-----------------------------------------------------------------------------
// Copyright (C) 2009 OutputLogic.com
// This source file may be used and distributed without restriction
// provided that this copyright statement is not removed from the file
// and that any derivative work contains the original copyright notice
// and the associated disclaimer.
//
// THIS SOURCE FILE IS PROVIDED "AS IS" AND WITHOUT ANY EXPRESS
// OR IMPLIED WARRANTIES, INCLUDING, WITHOUT LIMITATION, THE IMPLIED
// WARRANTIES OF MERCHANTIBILITY AND FITNESS FOR A PARTICULAR PURPOSE.
//-----------------------------------------------------------------------------
// CRC module for data[31:0] ,   crc[31:0]=1+x^1+x^2+x^4+x^5+x^7+x^8+x^10+x^11+x^12+x^16+x^22+x^23+x^26+x^32;
//-----------------------------------------------------------------------------

/* Allow valid byte valid for data_w == 16 */
module crc #(
	parameter DATA_W = 16,
	localparam KEEP_W = DATA_W/8,
	parameter LEN_W = $clog2(KEEP_W+1),
	parameter CRC_W = 32
)
(
  input               clk,
  input               valid_i,
  input  [LEN_W-1:0]  len_i,
  input               start_i,
  input  [DATA_W-1:0] data_i,
  output [CRC_W-1:0]  crc_o
);

  reg   [CRC_W-1:0] lfsr_q;
  logic [CRC_W-1:0] lfsr_next;
  logic [CRC_W-1:0] lfsr_next_arr[KEEP_W-1:0];
  logic [CRC_W-1:0] lfsr;

  assign crc_o = lfsr_q;
  assign lfsr = start_i ? {CRC_W{1'b1}} : lfsr_q;
if(DATA_W >= 8 ) begin

  assign lfsr_next_arr[0][0] = lfsr[24] ^ lfsr[30] ^ data_i[0] ^ data_i[6];
  assign lfsr_next_arr[0][1] = lfsr[24] ^ lfsr[25] ^ lfsr[30] ^ lfsr[31] ^ data_i[0] ^ data_i[1] ^ data_i[6] ^ data_i[7];
  assign lfsr_next_arr[0][2] = lfsr[24] ^ lfsr[25] ^ lfsr[26] ^ lfsr[30] ^ lfsr[31] ^ data_i[0] ^ data_i[1] ^ data_i[2] ^ data_i[6] ^ data_i[7];
  assign lfsr_next_arr[0][3] = lfsr[25] ^ lfsr[26] ^ lfsr[27] ^ lfsr[31] ^ data_i[1] ^ data_i[2] ^ data_i[3] ^ data_i[7];
  assign lfsr_next_arr[0][4] = lfsr[24] ^ lfsr[26] ^ lfsr[27] ^ lfsr[28] ^ lfsr[30] ^ data_i[0] ^ data_i[2] ^ data_i[3] ^ data_i[4] ^ data_i[6];
  assign lfsr_next_arr[0][5] = lfsr[24] ^ lfsr[25] ^ lfsr[27] ^ lfsr[28] ^ lfsr[29] ^ lfsr[30] ^ lfsr[31] ^ data_i[0] ^ data_i[1] ^ data_i[3] ^ data_i[4] ^ data_i[5] ^ data_i[6] ^ data_i[7];
  assign lfsr_next_arr[0][6] = lfsr[25] ^ lfsr[26] ^ lfsr[28] ^ lfsr[29] ^ lfsr[30] ^ lfsr[31] ^ data_i[1] ^ data_i[2] ^ data_i[4] ^ data_i[5] ^ data_i[6] ^ data_i[7];
  assign lfsr_next_arr[0][7] = lfsr[24] ^ lfsr[26] ^ lfsr[27] ^ lfsr[29] ^ lfsr[31] ^ data_i[0] ^ data_i[2] ^ data_i[3] ^ data_i[5] ^ data_i[7];
  assign lfsr_next_arr[0][8] = lfsr[0] ^ lfsr[24] ^ lfsr[25] ^ lfsr[27] ^ lfsr[28] ^ data_i[0] ^ data_i[1] ^ data_i[3] ^ data_i[4];
  assign lfsr_next_arr[0][9] = lfsr[1] ^ lfsr[25] ^ lfsr[26] ^ lfsr[28] ^ lfsr[29] ^ data_i[1] ^ data_i[2] ^ data_i[4] ^ data_i[5];
  assign lfsr_next_arr[0][10] = lfsr[2] ^ lfsr[24] ^ lfsr[26] ^ lfsr[27] ^ lfsr[29] ^ data_i[0] ^ data_i[2] ^ data_i[3] ^ data_i[5];
  assign lfsr_next_arr[0][11] = lfsr[3] ^ lfsr[24] ^ lfsr[25] ^ lfsr[27] ^ lfsr[28] ^ data_i[0] ^ data_i[1] ^ data_i[3] ^ data_i[4];
  assign lfsr_next_arr[0][12] = lfsr[4] ^ lfsr[24] ^ lfsr[25] ^ lfsr[26] ^ lfsr[28] ^ lfsr[29] ^ lfsr[30] ^ data_i[0] ^ data_i[1] ^ data_i[2] ^ data_i[4] ^ data_i[5] ^ data_i[6];
  assign lfsr_next_arr[0][13] = lfsr[5] ^ lfsr[25] ^ lfsr[26] ^ lfsr[27] ^ lfsr[29] ^ lfsr[30] ^ lfsr[31] ^ data_i[1] ^ data_i[2] ^ data_i[3] ^ data_i[5] ^ data_i[6] ^ data_i[7];
  assign lfsr_next_arr[0][14] = lfsr[6] ^ lfsr[26] ^ lfsr[27] ^ lfsr[28] ^ lfsr[30] ^ lfsr[31] ^ data_i[2] ^ data_i[3] ^ data_i[4] ^ data_i[6] ^ data_i[7];
  assign lfsr_next_arr[0][15] = lfsr[7] ^ lfsr[27] ^ lfsr[28] ^ lfsr[29] ^ lfsr[31] ^ data_i[3] ^ data_i[4] ^ data_i[5] ^ data_i[7];
  assign lfsr_next_arr[0][16] = lfsr[8] ^ lfsr[24] ^ lfsr[28] ^ lfsr[29] ^ data_i[0] ^ data_i[4] ^ data_i[5];
  assign lfsr_next_arr[0][17] = lfsr[9] ^ lfsr[25] ^ lfsr[29] ^ lfsr[30] ^ data_i[1] ^ data_i[5] ^ data_i[6];
  assign lfsr_next_arr[0][18] = lfsr[10] ^ lfsr[26] ^ lfsr[30] ^ lfsr[31] ^ data_i[2] ^ data_i[6] ^ data_i[7];
  assign lfsr_next_arr[0][19] = lfsr[11] ^ lfsr[27] ^ lfsr[31] ^ data_i[3] ^ data_i[7];
  assign lfsr_next_arr[0][20] = lfsr[12] ^ lfsr[28] ^ data_i[4];
  assign lfsr_next_arr[0][21] = lfsr[13] ^ lfsr[29] ^ data_i[5];
  assign lfsr_next_arr[0][22] = lfsr[14] ^ lfsr[24] ^ data_i[0];
  assign lfsr_next_arr[0][23] = lfsr[15] ^ lfsr[24] ^ lfsr[25] ^ lfsr[30] ^ data_i[0] ^ data_i[1] ^ data_i[6];
  assign lfsr_next_arr[0][24] = lfsr[16] ^ lfsr[25] ^ lfsr[26] ^ lfsr[31] ^ data_i[1] ^ data_i[2] ^ data_i[7];
  assign lfsr_next_arr[0][25] = lfsr[17] ^ lfsr[26] ^ lfsr[27] ^ data_i[2] ^ data_i[3];
  assign lfsr_next_arr[0][26] = lfsr[18] ^ lfsr[24] ^ lfsr[27] ^ lfsr[28] ^ lfsr[30] ^ data_i[0] ^ data_i[3] ^ data_i[4] ^ data_i[6];
  assign lfsr_next_arr[0][27] = lfsr[19] ^ lfsr[25] ^ lfsr[28] ^ lfsr[29] ^ lfsr[31] ^ data_i[1] ^ data_i[4] ^ data_i[5] ^ data_i[7];
  assign lfsr_next_arr[0][28] = lfsr[20] ^ lfsr[26] ^ lfsr[29] ^ lfsr[30] ^ data_i[2] ^ data_i[5] ^ data_i[6];
  assign lfsr_next_arr[0][29] = lfsr[21] ^ lfsr[27] ^ lfsr[30] ^ lfsr[31] ^ data_i[3] ^ data_i[6] ^ data_i[7];
  assign lfsr_next_arr[0][30] = lfsr[22] ^ lfsr[28] ^ lfsr[31] ^ data_i[4] ^ data_i[7];
  assign lfsr_next_arr[0][31] = lfsr[23] ^ lfsr[29] ^ data_i[5];

end 
if(DATA_W >= 16) begin

  assign  lfsr_next_arr[1][0] = lfsr[16] ^ lfsr[22] ^ lfsr[25] ^ lfsr[26] ^ lfsr[28] ^ data_i[0] ^ data_i[6] ^ data_i[9] ^ data_i[10] ^ data_i[12];
  assign  lfsr_next_arr[1][1] = lfsr[16] ^ lfsr[17] ^ lfsr[22] ^ lfsr[23] ^ lfsr[25] ^ lfsr[27] ^ lfsr[28] ^ lfsr[29] ^ data_i[0] ^ data_i[1] ^ data_i[6] ^ data_i[7] ^ data_i[9] ^ data_i[11] ^ data_i[12] ^ data_i[13];
  assign  lfsr_next_arr[1][2] = lfsr[16] ^ lfsr[17] ^ lfsr[18] ^ lfsr[22] ^ lfsr[23] ^ lfsr[24] ^ lfsr[25] ^ lfsr[29] ^ lfsr[30] ^ data_i[0] ^ data_i[1] ^ data_i[2] ^ data_i[6] ^ data_i[7] ^ data_i[8] ^ data_i[9] ^ data_i[13] ^ data_i[14];
  assign  lfsr_next_arr[1][3] = lfsr[17] ^ lfsr[18] ^ lfsr[19] ^ lfsr[23] ^ lfsr[24] ^ lfsr[25] ^ lfsr[26] ^ lfsr[30] ^ lfsr[31] ^ data_i[1] ^ data_i[2] ^ data_i[3] ^ data_i[7] ^ data_i[8] ^ data_i[9] ^ data_i[10] ^ data_i[14] ^ data_i[15];
  assign  lfsr_next_arr[1][4] = lfsr[16] ^ lfsr[18] ^ lfsr[19] ^ lfsr[20] ^ lfsr[22] ^ lfsr[24] ^ lfsr[27] ^ lfsr[28] ^ lfsr[31] ^ data_i[0] ^ data_i[2] ^ data_i[3] ^ data_i[4] ^ data_i[6] ^ data_i[8] ^ data_i[11] ^ data_i[12] ^ data_i[15];
  assign  lfsr_next_arr[1][5] = lfsr[16] ^ lfsr[17] ^ lfsr[19] ^ lfsr[20] ^ lfsr[21] ^ lfsr[22] ^ lfsr[23] ^ lfsr[26] ^ lfsr[29] ^ data_i[0] ^ data_i[1] ^ data_i[3] ^ data_i[4] ^ data_i[5] ^ data_i[6] ^ data_i[7] ^ data_i[10] ^ data_i[13];
  assign  lfsr_next_arr[1][6] = lfsr[17] ^ lfsr[18] ^ lfsr[20] ^ lfsr[21] ^ lfsr[22] ^ lfsr[23] ^ lfsr[24] ^ lfsr[27] ^ lfsr[30] ^ data_i[1] ^ data_i[2] ^ data_i[4] ^ data_i[5] ^ data_i[6] ^ data_i[7] ^ data_i[8] ^ data_i[11] ^ data_i[14];
  assign  lfsr_next_arr[1][7] = lfsr[16] ^ lfsr[18] ^ lfsr[19] ^ lfsr[21] ^ lfsr[23] ^ lfsr[24] ^ lfsr[26] ^ lfsr[31] ^ data_i[0] ^ data_i[2] ^ data_i[3] ^ data_i[5] ^ data_i[7] ^ data_i[8] ^ data_i[10] ^ data_i[15];
  assign  lfsr_next_arr[1][8] = lfsr[16] ^ lfsr[17] ^ lfsr[19] ^ lfsr[20] ^ lfsr[24] ^ lfsr[26] ^ lfsr[27] ^ lfsr[28] ^ data_i[0] ^ data_i[1] ^ data_i[3] ^ data_i[4] ^ data_i[8] ^ data_i[10] ^ data_i[11] ^ data_i[12];
  assign  lfsr_next_arr[1][9] = lfsr[17] ^ lfsr[18] ^ lfsr[20] ^ lfsr[21] ^ lfsr[25] ^ lfsr[27] ^ lfsr[28] ^ lfsr[29] ^ data_i[1] ^ data_i[2] ^ data_i[4] ^ data_i[5] ^ data_i[9] ^ data_i[11] ^ data_i[12] ^ data_i[13];
  assign  lfsr_next_arr[1][10] = lfsr[16] ^ lfsr[18] ^ lfsr[19] ^ lfsr[21] ^ lfsr[25] ^ lfsr[29] ^ lfsr[30] ^ data_i[0] ^ data_i[2] ^ data_i[3] ^ data_i[5] ^ data_i[9] ^ data_i[13] ^ data_i[14];
  assign  lfsr_next_arr[1][11] = lfsr[16] ^ lfsr[17] ^ lfsr[19] ^ lfsr[20] ^ lfsr[25] ^ lfsr[28] ^ lfsr[30] ^ lfsr[31] ^ data_i[0] ^ data_i[1] ^ data_i[3] ^ data_i[4] ^ data_i[9] ^ data_i[12] ^ data_i[14] ^ data_i[15];
  assign  lfsr_next_arr[1][12] = lfsr[16] ^ lfsr[17] ^ lfsr[18] ^ lfsr[20] ^ lfsr[21] ^ lfsr[22] ^ lfsr[25] ^ lfsr[28] ^ lfsr[29] ^ lfsr[31] ^ data_i[0] ^ data_i[1] ^ data_i[2] ^ data_i[4] ^ data_i[5] ^ data_i[6] ^ data_i[9] ^ data_i[12] ^ data_i[13] ^ data_i[15];
  assign  lfsr_next_arr[1][13] = lfsr[17] ^ lfsr[18] ^ lfsr[19] ^ lfsr[21] ^ lfsr[22] ^ lfsr[23] ^ lfsr[26] ^ lfsr[29] ^ lfsr[30] ^ data_i[1] ^ data_i[2] ^ data_i[3] ^ data_i[5] ^ data_i[6] ^ data_i[7] ^ data_i[10] ^ data_i[13] ^ data_i[14];
  assign  lfsr_next_arr[1][14] = lfsr[18] ^ lfsr[19] ^ lfsr[20] ^ lfsr[22] ^ lfsr[23] ^ lfsr[24] ^ lfsr[27] ^ lfsr[30] ^ lfsr[31] ^ data_i[2] ^ data_i[3] ^ data_i[4] ^ data_i[6] ^ data_i[7] ^ data_i[8] ^ data_i[11] ^ data_i[14] ^ data_i[15];
  assign  lfsr_next_arr[1][15] = lfsr[19] ^ lfsr[20] ^ lfsr[21] ^ lfsr[23] ^ lfsr[24] ^ lfsr[25] ^ lfsr[28] ^ lfsr[31] ^ data_i[3] ^ data_i[4] ^ data_i[5] ^ data_i[7] ^ data_i[8] ^ data_i[9] ^ data_i[12] ^ data_i[15];
  assign  lfsr_next_arr[1][16] = lfsr[0] ^ lfsr[16] ^ lfsr[20] ^ lfsr[21] ^ lfsr[24] ^ lfsr[28] ^ lfsr[29] ^ data_i[0] ^ data_i[4] ^ data_i[5] ^ data_i[8] ^ data_i[12] ^ data_i[13];
  assign  lfsr_next_arr[1][17] = lfsr[1] ^ lfsr[17] ^ lfsr[21] ^ lfsr[22] ^ lfsr[25] ^ lfsr[29] ^ lfsr[30] ^ data_i[1] ^ data_i[5] ^ data_i[6] ^ data_i[9] ^ data_i[13] ^ data_i[14];
  assign  lfsr_next_arr[1][18] = lfsr[2] ^ lfsr[18] ^ lfsr[22] ^ lfsr[23] ^ lfsr[26] ^ lfsr[30] ^ lfsr[31] ^ data_i[2] ^ data_i[6] ^ data_i[7] ^ data_i[10] ^ data_i[14] ^ data_i[15];
  assign  lfsr_next_arr[1][19] = lfsr[3] ^ lfsr[19] ^ lfsr[23] ^ lfsr[24] ^ lfsr[27] ^ lfsr[31] ^ data_i[3] ^ data_i[7] ^ data_i[8] ^ data_i[11] ^ data_i[15];
  assign  lfsr_next_arr[1][20] = lfsr[4] ^ lfsr[20] ^ lfsr[24] ^ lfsr[25] ^ lfsr[28] ^ data_i[4] ^ data_i[8] ^ data_i[9] ^ data_i[12];
  assign  lfsr_next_arr[1][21] = lfsr[5] ^ lfsr[21] ^ lfsr[25] ^ lfsr[26] ^ lfsr[29] ^ data_i[5] ^ data_i[9] ^ data_i[10] ^ data_i[13];
  assign  lfsr_next_arr[1][22] = lfsr[6] ^ lfsr[16] ^ lfsr[25] ^ lfsr[27] ^ lfsr[28] ^ lfsr[30] ^ data_i[0] ^ data_i[9] ^ data_i[11] ^ data_i[12] ^ data_i[14];
  assign  lfsr_next_arr[1][23] = lfsr[7] ^ lfsr[16] ^ lfsr[17] ^ lfsr[22] ^ lfsr[25] ^ lfsr[29] ^ lfsr[31] ^ data_i[0] ^ data_i[1] ^ data_i[6] ^ data_i[9] ^ data_i[13] ^ data_i[15];
  assign  lfsr_next_arr[1][24] = lfsr[8] ^ lfsr[17] ^ lfsr[18] ^ lfsr[23] ^ lfsr[26] ^ lfsr[30] ^ data_i[1] ^ data_i[2] ^ data_i[7] ^ data_i[10] ^ data_i[14];
  assign  lfsr_next_arr[1][25] = lfsr[9] ^ lfsr[18] ^ lfsr[19] ^ lfsr[24] ^ lfsr[27] ^ lfsr[31] ^ data_i[2] ^ data_i[3] ^ data_i[8] ^ data_i[11] ^ data_i[15];
  assign  lfsr_next_arr[1][26] = lfsr[10] ^ lfsr[16] ^ lfsr[19] ^ lfsr[20] ^ lfsr[22] ^ lfsr[26] ^ data_i[0] ^ data_i[3] ^ data_i[4] ^ data_i[6] ^ data_i[10];
  assign  lfsr_next_arr[1][27] = lfsr[11] ^ lfsr[17] ^ lfsr[20] ^ lfsr[21] ^ lfsr[23] ^ lfsr[27] ^ data_i[1] ^ data_i[4] ^ data_i[5] ^ data_i[7] ^ data_i[11];
  assign  lfsr_next_arr[1][28] = lfsr[12] ^ lfsr[18] ^ lfsr[21] ^ lfsr[22] ^ lfsr[24] ^ lfsr[28] ^ data_i[2] ^ data_i[5] ^ data_i[6] ^ data_i[8] ^ data_i[12];
  assign  lfsr_next_arr[1][29] = lfsr[13] ^ lfsr[19] ^ lfsr[22] ^ lfsr[23] ^ lfsr[25] ^ lfsr[29] ^ data_i[3] ^ data_i[6] ^ data_i[7] ^ data_i[9] ^ data_i[13];
  assign  lfsr_next_arr[1][30] = lfsr[14] ^ lfsr[20] ^ lfsr[23] ^ lfsr[24] ^ lfsr[26] ^ lfsr[30] ^ data_i[4] ^ data_i[7] ^ data_i[8] ^ data_i[10] ^ data_i[14];
  assign  lfsr_next_arr[1][31] = lfsr[15] ^ lfsr[21] ^ lfsr[24] ^ lfsr[25] ^ lfsr[27] ^ lfsr[31] ^ data_i[5] ^ data_i[8] ^ data_i[9] ^ data_i[11] ^ data_i[15];

end 
if(DATA_W == 32) begin

   assign lfsr_next_arr[3][0] = lfsr[0] ^ lfsr[6] ^ lfsr[9] ^ lfsr[10] ^ lfsr[12] ^ lfsr[16] ^ lfsr[24] ^ lfsr[25] ^ lfsr[26] ^ lfsr[28] ^ lfsr[29] ^ lfsr[30] ^ lfsr[31] ^ data_i[0] ^ data_i[6] ^ data_i[9] ^ data_i[10] ^ data_i[12] ^ data_i[16] ^ data_i[24] ^ data_i[25] ^ data_i[26] ^ data_i[28] ^ data_i[29] ^ data_i[30] ^ data_i[31];
   assign lfsr_next_arr[3][1] = lfsr[0] ^ lfsr[1] ^ lfsr[6] ^ lfsr[7] ^ lfsr[9] ^ lfsr[11] ^ lfsr[12] ^ lfsr[13] ^ lfsr[16] ^ lfsr[17] ^ lfsr[24] ^ lfsr[27] ^ lfsr[28] ^ data_i[0] ^ data_i[1] ^ data_i[6] ^ data_i[7] ^ data_i[9] ^ data_i[11] ^ data_i[12] ^ data_i[13] ^ data_i[16] ^ data_i[17] ^ data_i[24] ^ data_i[27] ^ data_i[28];
   assign lfsr_next_arr[3][2] = lfsr[0] ^ lfsr[1] ^ lfsr[2] ^ lfsr[6] ^ lfsr[7] ^ lfsr[8] ^ lfsr[9] ^ lfsr[13] ^ lfsr[14] ^ lfsr[16] ^ lfsr[17] ^ lfsr[18] ^ lfsr[24] ^ lfsr[26] ^ lfsr[30] ^ lfsr[31] ^ data_i[0] ^ data_i[1] ^ data_i[2] ^ data_i[6] ^ data_i[7] ^ data_i[8] ^ data_i[9] ^ data_i[13] ^ data_i[14] ^ data_i[16] ^ data_i[17] ^ data_i[18] ^ data_i[24] ^ data_i[26] ^ data_i[30] ^ data_i[31];
   assign lfsr_next_arr[3][3] = lfsr[1] ^ lfsr[2] ^ lfsr[3] ^ lfsr[7] ^ lfsr[8] ^ lfsr[9] ^ lfsr[10] ^ lfsr[14] ^ lfsr[15] ^ lfsr[17] ^ lfsr[18] ^ lfsr[19] ^ lfsr[25] ^ lfsr[27] ^ lfsr[31] ^ data_i[1] ^ data_i[2] ^ data_i[3] ^ data_i[7] ^ data_i[8] ^ data_i[9] ^ data_i[10] ^ data_i[14] ^ data_i[15] ^ data_i[17] ^ data_i[18] ^ data_i[19] ^ data_i[25] ^ data_i[27] ^ data_i[31];
   assign lfsr_next_arr[3][4] = lfsr[0] ^ lfsr[2] ^ lfsr[3] ^ lfsr[4] ^ lfsr[6] ^ lfsr[8] ^ lfsr[11] ^ lfsr[12] ^ lfsr[15] ^ lfsr[18] ^ lfsr[19] ^ lfsr[20] ^ lfsr[24] ^ lfsr[25] ^ lfsr[29] ^ lfsr[30] ^ lfsr[31] ^ data_i[0] ^ data_i[2] ^ data_i[3] ^ data_i[4] ^ data_i[6] ^ data_i[8] ^ data_i[11] ^ data_i[12] ^ data_i[15] ^ data_i[18] ^ data_i[19] ^ data_i[20] ^ data_i[24] ^ data_i[25] ^ data_i[29] ^ data_i[30] ^ data_i[31];
   assign lfsr_next_arr[3][5] = lfsr[0] ^ lfsr[1] ^ lfsr[3] ^ lfsr[4] ^ lfsr[5] ^ lfsr[6] ^ lfsr[7] ^ lfsr[10] ^ lfsr[13] ^ lfsr[19] ^ lfsr[20] ^ lfsr[21] ^ lfsr[24] ^ lfsr[28] ^ lfsr[29] ^ data_i[0] ^ data_i[1] ^ data_i[3] ^ data_i[4] ^ data_i[5] ^ data_i[6] ^ data_i[7] ^ data_i[10] ^ data_i[13] ^ data_i[19] ^ data_i[20] ^ data_i[21] ^ data_i[24] ^ data_i[28] ^ data_i[29];
   assign lfsr_next_arr[3][6] = lfsr[1] ^ lfsr[2] ^ lfsr[4] ^ lfsr[5] ^ lfsr[6] ^ lfsr[7] ^ lfsr[8] ^ lfsr[11] ^ lfsr[14] ^ lfsr[20] ^ lfsr[21] ^ lfsr[22] ^ lfsr[25] ^ lfsr[29] ^ lfsr[30] ^ data_i[1] ^ data_i[2] ^ data_i[4] ^ data_i[5] ^ data_i[6] ^ data_i[7] ^ data_i[8] ^ data_i[11] ^ data_i[14] ^ data_i[20] ^ data_i[21] ^ data_i[22] ^ data_i[25] ^ data_i[29] ^ data_i[30];
   assign lfsr_next_arr[3][7] = lfsr[0] ^ lfsr[2] ^ lfsr[3] ^ lfsr[5] ^ lfsr[7] ^ lfsr[8] ^ lfsr[10] ^ lfsr[15] ^ lfsr[16] ^ lfsr[21] ^ lfsr[22] ^ lfsr[23] ^ lfsr[24] ^ lfsr[25] ^ lfsr[28] ^ lfsr[29] ^ data_i[0] ^ data_i[2] ^ data_i[3] ^ data_i[5] ^ data_i[7] ^ data_i[8] ^ data_i[10] ^ data_i[15] ^ data_i[16] ^ data_i[21] ^ data_i[22] ^ data_i[23] ^ data_i[24] ^ data_i[25] ^ data_i[28] ^ data_i[29];
   assign lfsr_next_arr[3][8] = lfsr[0] ^ lfsr[1] ^ lfsr[3] ^ lfsr[4] ^ lfsr[8] ^ lfsr[10] ^ lfsr[11] ^ lfsr[12] ^ lfsr[17] ^ lfsr[22] ^ lfsr[23] ^ lfsr[28] ^ lfsr[31] ^ data_i[0] ^ data_i[1] ^ data_i[3] ^ data_i[4] ^ data_i[8] ^ data_i[10] ^ data_i[11] ^ data_i[12] ^ data_i[17] ^ data_i[22] ^ data_i[23] ^ data_i[28] ^ data_i[31];
   assign lfsr_next_arr[3][9] = lfsr[1] ^ lfsr[2] ^ lfsr[4] ^ lfsr[5] ^ lfsr[9] ^ lfsr[11] ^ lfsr[12] ^ lfsr[13] ^ lfsr[18] ^ lfsr[23] ^ lfsr[24] ^ lfsr[29] ^ data_i[1] ^ data_i[2] ^ data_i[4] ^ data_i[5] ^ data_i[9] ^ data_i[11] ^ data_i[12] ^ data_i[13] ^ data_i[18] ^ data_i[23] ^ data_i[24] ^ data_i[29];
   assign lfsr_next_arr[3][10] = lfsr[0] ^ lfsr[2] ^ lfsr[3] ^ lfsr[5] ^ lfsr[9] ^ lfsr[13] ^ lfsr[14] ^ lfsr[16] ^ lfsr[19] ^ lfsr[26] ^ lfsr[28] ^ lfsr[29] ^ lfsr[31] ^ data_i[0] ^ data_i[2] ^ data_i[3] ^ data_i[5] ^ data_i[9] ^ data_i[13] ^ data_i[14] ^ data_i[16] ^ data_i[19] ^ data_i[26] ^ data_i[28] ^ data_i[29] ^ data_i[31];
   assign lfsr_next_arr[3][11] = lfsr[0] ^ lfsr[1] ^ lfsr[3] ^ lfsr[4] ^ lfsr[9] ^ lfsr[12] ^ lfsr[14] ^ lfsr[15] ^ lfsr[16] ^ lfsr[17] ^ lfsr[20] ^ lfsr[24] ^ lfsr[25] ^ lfsr[26] ^ lfsr[27] ^ lfsr[28] ^ lfsr[31] ^ data_i[0] ^ data_i[1] ^ data_i[3] ^ data_i[4] ^ data_i[9] ^ data_i[12] ^ data_i[14] ^ data_i[15] ^ data_i[16] ^ data_i[17] ^ data_i[20] ^ data_i[24] ^ data_i[25] ^ data_i[26] ^ data_i[27] ^ data_i[28] ^ data_i[31];
   assign lfsr_next_arr[3][12] = lfsr[0] ^ lfsr[1] ^ lfsr[2] ^ lfsr[4] ^ lfsr[5] ^ lfsr[6] ^ lfsr[9] ^ lfsr[12] ^ lfsr[13] ^ lfsr[15] ^ lfsr[17] ^ lfsr[18] ^ lfsr[21] ^ lfsr[24] ^ lfsr[27] ^ lfsr[30] ^ lfsr[31] ^ data_i[0] ^ data_i[1] ^ data_i[2] ^ data_i[4] ^ data_i[5] ^ data_i[6] ^ data_i[9] ^ data_i[12] ^ data_i[13] ^ data_i[15] ^ data_i[17] ^ data_i[18] ^ data_i[21] ^ data_i[24] ^ data_i[27] ^ data_i[30] ^ data_i[31];
   assign lfsr_next_arr[3][13] = lfsr[1] ^ lfsr[2] ^ lfsr[3] ^ lfsr[5] ^ lfsr[6] ^ lfsr[7] ^ lfsr[10] ^ lfsr[13] ^ lfsr[14] ^ lfsr[16] ^ lfsr[18] ^ lfsr[19] ^ lfsr[22] ^ lfsr[25] ^ lfsr[28] ^ lfsr[31] ^ data_i[1] ^ data_i[2] ^ data_i[3] ^ data_i[5] ^ data_i[6] ^ data_i[7] ^ data_i[10] ^ data_i[13] ^ data_i[14] ^ data_i[16] ^ data_i[18] ^ data_i[19] ^ data_i[22] ^ data_i[25] ^ data_i[28] ^ data_i[31];
   assign lfsr_next_arr[3][14] = lfsr[2] ^ lfsr[3] ^ lfsr[4] ^ lfsr[6] ^ lfsr[7] ^ lfsr[8] ^ lfsr[11] ^ lfsr[14] ^ lfsr[15] ^ lfsr[17] ^ lfsr[19] ^ lfsr[20] ^ lfsr[23] ^ lfsr[26] ^ lfsr[29] ^ data_i[2] ^ data_i[3] ^ data_i[4] ^ data_i[6] ^ data_i[7] ^ data_i[8] ^ data_i[11] ^ data_i[14] ^ data_i[15] ^ data_i[17] ^ data_i[19] ^ data_i[20] ^ data_i[23] ^ data_i[26] ^ data_i[29];
   assign lfsr_next_arr[3][15] = lfsr[3] ^ lfsr[4] ^ lfsr[5] ^ lfsr[7] ^ lfsr[8] ^ lfsr[9] ^ lfsr[12] ^ lfsr[15] ^ lfsr[16] ^ lfsr[18] ^ lfsr[20] ^ lfsr[21] ^ lfsr[24] ^ lfsr[27] ^ lfsr[30] ^ data_i[3] ^ data_i[4] ^ data_i[5] ^ data_i[7] ^ data_i[8] ^ data_i[9] ^ data_i[12] ^ data_i[15] ^ data_i[16] ^ data_i[18] ^ data_i[20] ^ data_i[21] ^ data_i[24] ^ data_i[27] ^ data_i[30];
   assign lfsr_next_arr[3][16] = lfsr[0] ^ lfsr[4] ^ lfsr[5] ^ lfsr[8] ^ lfsr[12] ^ lfsr[13] ^ lfsr[17] ^ lfsr[19] ^ lfsr[21] ^ lfsr[22] ^ lfsr[24] ^ lfsr[26] ^ lfsr[29] ^ lfsr[30] ^ data_i[0] ^ data_i[4] ^ data_i[5] ^ data_i[8] ^ data_i[12] ^ data_i[13] ^ data_i[17] ^ data_i[19] ^ data_i[21] ^ data_i[22] ^ data_i[24] ^ data_i[26] ^ data_i[29] ^ data_i[30];
   assign lfsr_next_arr[3][17] = lfsr[1] ^ lfsr[5] ^ lfsr[6] ^ lfsr[9] ^ lfsr[13] ^ lfsr[14] ^ lfsr[18] ^ lfsr[20] ^ lfsr[22] ^ lfsr[23] ^ lfsr[25] ^ lfsr[27] ^ lfsr[30] ^ lfsr[31] ^ data_i[1] ^ data_i[5] ^ data_i[6] ^ data_i[9] ^ data_i[13] ^ data_i[14] ^ data_i[18] ^ data_i[20] ^ data_i[22] ^ data_i[23] ^ data_i[25] ^ data_i[27] ^ data_i[30] ^ data_i[31];
   assign lfsr_next_arr[3][18] = lfsr[2] ^ lfsr[6] ^ lfsr[7] ^ lfsr[10] ^ lfsr[14] ^ lfsr[15] ^ lfsr[19] ^ lfsr[21] ^ lfsr[23] ^ lfsr[24] ^ lfsr[26] ^ lfsr[28] ^ lfsr[31] ^ data_i[2] ^ data_i[6] ^ data_i[7] ^ data_i[10] ^ data_i[14] ^ data_i[15] ^ data_i[19] ^ data_i[21] ^ data_i[23] ^ data_i[24] ^ data_i[26] ^ data_i[28] ^ data_i[31];
   assign lfsr_next_arr[3][19] = lfsr[3] ^ lfsr[7] ^ lfsr[8] ^ lfsr[11] ^ lfsr[15] ^ lfsr[16] ^ lfsr[20] ^ lfsr[22] ^ lfsr[24] ^ lfsr[25] ^ lfsr[27] ^ lfsr[29] ^ data_i[3] ^ data_i[7] ^ data_i[8] ^ data_i[11] ^ data_i[15] ^ data_i[16] ^ data_i[20] ^ data_i[22] ^ data_i[24] ^ data_i[25] ^ data_i[27] ^ data_i[29];
   assign lfsr_next_arr[3][20] = lfsr[4] ^ lfsr[8] ^ lfsr[9] ^ lfsr[12] ^ lfsr[16] ^ lfsr[17] ^ lfsr[21] ^ lfsr[23] ^ lfsr[25] ^ lfsr[26] ^ lfsr[28] ^ lfsr[30] ^ data_i[4] ^ data_i[8] ^ data_i[9] ^ data_i[12] ^ data_i[16] ^ data_i[17] ^ data_i[21] ^ data_i[23] ^ data_i[25] ^ data_i[26] ^ data_i[28] ^ data_i[30];
   assign lfsr_next_arr[3][21] = lfsr[5] ^ lfsr[9] ^ lfsr[10] ^ lfsr[13] ^ lfsr[17] ^ lfsr[18] ^ lfsr[22] ^ lfsr[24] ^ lfsr[26] ^ lfsr[27] ^ lfsr[29] ^ lfsr[31] ^ data_i[5] ^ data_i[9] ^ data_i[10] ^ data_i[13] ^ data_i[17] ^ data_i[18] ^ data_i[22] ^ data_i[24] ^ data_i[26] ^ data_i[27] ^ data_i[29] ^ data_i[31];
   assign lfsr_next_arr[3][22] = lfsr[0] ^ lfsr[9] ^ lfsr[11] ^ lfsr[12] ^ lfsr[14] ^ lfsr[16] ^ lfsr[18] ^ lfsr[19] ^ lfsr[23] ^ lfsr[24] ^ lfsr[26] ^ lfsr[27] ^ lfsr[29] ^ lfsr[31] ^ data_i[0] ^ data_i[9] ^ data_i[11] ^ data_i[12] ^ data_i[14] ^ data_i[16] ^ data_i[18] ^ data_i[19] ^ data_i[23] ^ data_i[24] ^ data_i[26] ^ data_i[27] ^ data_i[29] ^ data_i[31];
   assign lfsr_next_arr[3][23] = lfsr[0] ^ lfsr[1] ^ lfsr[6] ^ lfsr[9] ^ lfsr[13] ^ lfsr[15] ^ lfsr[16] ^ lfsr[17] ^ lfsr[19] ^ lfsr[20] ^ lfsr[26] ^ lfsr[27] ^ lfsr[29] ^ lfsr[31] ^ data_i[0] ^ data_i[1] ^ data_i[6] ^ data_i[9] ^ data_i[13] ^ data_i[15] ^ data_i[16] ^ data_i[17] ^ data_i[19] ^ data_i[20] ^ data_i[26] ^ data_i[27] ^ data_i[29] ^ data_i[31];
   assign lfsr_next_arr[3][24] = lfsr[1] ^ lfsr[2] ^ lfsr[7] ^ lfsr[10] ^ lfsr[14] ^ lfsr[16] ^ lfsr[17] ^ lfsr[18] ^ lfsr[20] ^ lfsr[21] ^ lfsr[27] ^ lfsr[28] ^ lfsr[30] ^ data_i[1] ^ data_i[2] ^ data_i[7] ^ data_i[10] ^ data_i[14] ^ data_i[16] ^ data_i[17] ^ data_i[18] ^ data_i[20] ^ data_i[21] ^ data_i[27] ^ data_i[28] ^ data_i[30];
   assign lfsr_next_arr[3][25] = lfsr[2] ^ lfsr[3] ^ lfsr[8] ^ lfsr[11] ^ lfsr[15] ^ lfsr[17] ^ lfsr[18] ^ lfsr[19] ^ lfsr[21] ^ lfsr[22] ^ lfsr[28] ^ lfsr[29] ^ lfsr[31] ^ data_i[2] ^ data_i[3] ^ data_i[8] ^ data_i[11] ^ data_i[15] ^ data_i[17] ^ data_i[18] ^ data_i[19] ^ data_i[21] ^ data_i[22] ^ data_i[28] ^ data_i[29] ^ data_i[31];
   assign lfsr_next_arr[3][26] = lfsr[0] ^ lfsr[3] ^ lfsr[4] ^ lfsr[6] ^ lfsr[10] ^ lfsr[18] ^ lfsr[19] ^ lfsr[20] ^ lfsr[22] ^ lfsr[23] ^ lfsr[24] ^ lfsr[25] ^ lfsr[26] ^ lfsr[28] ^ lfsr[31] ^ data_i[0] ^ data_i[3] ^ data_i[4] ^ data_i[6] ^ data_i[10] ^ data_i[18] ^ data_i[19] ^ data_i[20] ^ data_i[22] ^ data_i[23] ^ data_i[24] ^ data_i[25] ^ data_i[26] ^ data_i[28] ^ data_i[31];
   assign lfsr_next_arr[3][27] = lfsr[1] ^ lfsr[4] ^ lfsr[5] ^ lfsr[7] ^ lfsr[11] ^ lfsr[19] ^ lfsr[20] ^ lfsr[21] ^ lfsr[23] ^ lfsr[24] ^ lfsr[25] ^ lfsr[26] ^ lfsr[27] ^ lfsr[29] ^ data_i[1] ^ data_i[4] ^ data_i[5] ^ data_i[7] ^ data_i[11] ^ data_i[19] ^ data_i[20] ^ data_i[21] ^ data_i[23] ^ data_i[24] ^ data_i[25] ^ data_i[26] ^ data_i[27] ^ data_i[29];
   assign lfsr_next_arr[3][28] = lfsr[2] ^ lfsr[5] ^ lfsr[6] ^ lfsr[8] ^ lfsr[12] ^ lfsr[20] ^ lfsr[21] ^ lfsr[22] ^ lfsr[24] ^ lfsr[25] ^ lfsr[26] ^ lfsr[27] ^ lfsr[28] ^ lfsr[30] ^ data_i[2] ^ data_i[5] ^ data_i[6] ^ data_i[8] ^ data_i[12] ^ data_i[20] ^ data_i[21] ^ data_i[22] ^ data_i[24] ^ data_i[25] ^ data_i[26] ^ data_i[27] ^ data_i[28] ^ data_i[30];
   assign lfsr_next_arr[3][29] = lfsr[3] ^ lfsr[6] ^ lfsr[7] ^ lfsr[9] ^ lfsr[13] ^ lfsr[21] ^ lfsr[22] ^ lfsr[23] ^ lfsr[25] ^ lfsr[26] ^ lfsr[27] ^ lfsr[28] ^ lfsr[29] ^ lfsr[31] ^ data_i[3] ^ data_i[6] ^ data_i[7] ^ data_i[9] ^ data_i[13] ^ data_i[21] ^ data_i[22] ^ data_i[23] ^ data_i[25] ^ data_i[26] ^ data_i[27] ^ data_i[28] ^ data_i[29] ^ data_i[31];
   assign lfsr_next_arr[3][30] = lfsr[4] ^ lfsr[7] ^ lfsr[8] ^ lfsr[10] ^ lfsr[14] ^ lfsr[22] ^ lfsr[23] ^ lfsr[24] ^ lfsr[26] ^ lfsr[27] ^ lfsr[28] ^ lfsr[29] ^ lfsr[30] ^ data_i[4] ^ data_i[7] ^ data_i[8] ^ data_i[10] ^ data_i[14] ^ data_i[22] ^ data_i[23] ^ data_i[24] ^ data_i[26] ^ data_i[27] ^ data_i[28] ^ data_i[29] ^ data_i[30];
   assign lfsr_next_arr[3][31] = lfsr[5] ^ lfsr[8] ^ lfsr[9] ^ lfsr[11] ^ lfsr[15] ^ lfsr[23] ^ lfsr[24] ^ lfsr[25] ^ lfsr[27] ^ lfsr[28] ^ lfsr[29] ^ lfsr[30] ^ lfsr[31] ^ data_i[5] ^ data_i[8] ^ data_i[9] ^ data_i[11] ^ data_i[15] ^ data_i[23] ^ data_i[24] ^ data_i[25] ^ data_i[27] ^ data_i[28] ^ data_i[29] ^ data_i[30] ^ data_i[31];

end 
if ( DATA_W == 64 ) begin

	assign lfsr_next_arr[7][0] = lfsr[0] ^ lfsr[2] ^ lfsr[5] ^ lfsr[12] ^ lfsr[13] ^ lfsr[15] ^ lfsr[16] ^ lfsr[18] ^ lfsr[21] ^ lfsr[22] ^ lfsr[23] ^ lfsr[26] ^ lfsr[28] ^ lfsr[29] ^ lfsr[31] ^ data_i[0] ^ data_i[6] ^ data_i[9] ^ data_i[10] ^ data_i[12] ^ data_i[16] ^ data_i[24] ^ data_i[25] ^ data_i[26] ^ data_i[28] ^ data_i[29] ^ data_i[30] ^ data_i[31] ^ data_i[32] ^ data_i[34] ^ data_i[37] ^ data_i[44] ^ data_i[45] ^ data_i[47] ^ data_i[48] ^ data_i[50] ^ data_i[53] ^ data_i[54] ^ data_i[55] ^ data_i[58] ^ data_i[60] ^ data_i[61] ^ data_i[63];
    assign lfsr_next_arr[7][1] = lfsr[1] ^ lfsr[2] ^ lfsr[3] ^ lfsr[5] ^ lfsr[6] ^ lfsr[12] ^ lfsr[14] ^ lfsr[15] ^ lfsr[17] ^ lfsr[18] ^ lfsr[19] ^ lfsr[21] ^ lfsr[24] ^ lfsr[26] ^ lfsr[27] ^ lfsr[28] ^ lfsr[30] ^ lfsr[31] ^ data_i[0] ^ data_i[1] ^ data_i[6] ^ data_i[7] ^ data_i[9] ^ data_i[11] ^ data_i[12] ^ data_i[13] ^ data_i[16] ^ data_i[17] ^ data_i[24] ^ data_i[27] ^ data_i[28] ^ data_i[33] ^ data_i[34] ^ data_i[35] ^ data_i[37] ^ data_i[38] ^ data_i[44] ^ data_i[46] ^ data_i[47] ^ data_i[49] ^ data_i[50] ^ data_i[51] ^ data_i[53] ^ data_i[56] ^ data_i[58] ^ data_i[59] ^ data_i[60] ^ data_i[62] ^ data_i[63];
    assign lfsr_next_arr[7][2] = lfsr[0] ^ lfsr[3] ^ lfsr[4] ^ lfsr[5] ^ lfsr[6] ^ lfsr[7] ^ lfsr[12] ^ lfsr[19] ^ lfsr[20] ^ lfsr[21] ^ lfsr[23] ^ lfsr[25] ^ lfsr[26] ^ lfsr[27] ^ data_i[0] ^ data_i[1] ^ data_i[2] ^ data_i[6] ^ data_i[7] ^ data_i[8] ^ data_i[9] ^ data_i[13] ^ data_i[14] ^ data_i[16] ^ data_i[17] ^ data_i[18] ^ data_i[24] ^ data_i[26] ^ data_i[30] ^ data_i[31] ^ data_i[32] ^ data_i[35] ^ data_i[36] ^ data_i[37] ^ data_i[38] ^ data_i[39] ^ data_i[44] ^ data_i[51] ^ data_i[52] ^ data_i[53] ^ data_i[55] ^ data_i[57] ^ data_i[58] ^ data_i[59];
    assign lfsr_next_arr[7][3] = lfsr[0] ^ lfsr[1] ^ lfsr[4] ^ lfsr[5] ^ lfsr[6] ^ lfsr[7] ^ lfsr[8] ^ lfsr[13] ^ lfsr[20] ^ lfsr[21] ^ lfsr[22] ^ lfsr[24] ^ lfsr[26] ^ lfsr[27] ^ lfsr[28] ^ data_i[1] ^ data_i[2] ^ data_i[3] ^ data_i[7] ^ data_i[8] ^ data_i[9] ^ data_i[10] ^ data_i[14] ^ data_i[15] ^ data_i[17] ^ data_i[18] ^ data_i[19] ^ data_i[25] ^ data_i[27] ^ data_i[31] ^ data_i[32] ^ data_i[33] ^ data_i[36] ^ data_i[37] ^ data_i[38] ^ data_i[39] ^ data_i[40] ^ data_i[45] ^ data_i[52] ^ data_i[53] ^ data_i[54] ^ data_i[56] ^ data_i[58] ^ data_i[59] ^ data_i[60];
    assign lfsr_next_arr[7][4] = lfsr[1] ^ lfsr[6] ^ lfsr[7] ^ lfsr[8] ^ lfsr[9] ^ lfsr[12] ^ lfsr[13] ^ lfsr[14] ^ lfsr[15] ^ lfsr[16] ^ lfsr[18] ^ lfsr[25] ^ lfsr[26] ^ lfsr[27] ^ lfsr[31] ^ data_i[0] ^ data_i[2] ^ data_i[3] ^ data_i[4] ^ data_i[6] ^ data_i[8] ^ data_i[11] ^ data_i[12] ^ data_i[15] ^ data_i[18] ^ data_i[19] ^ data_i[20] ^ data_i[24] ^ data_i[25] ^ data_i[29] ^ data_i[30] ^ data_i[31] ^ data_i[33] ^ data_i[38] ^ data_i[39] ^ data_i[40] ^ data_i[41] ^ data_i[44] ^ data_i[45] ^ data_i[46] ^ data_i[47] ^ data_i[48] ^ data_i[50] ^ data_i[57] ^ data_i[58] ^ data_i[59] ^ data_i[63];
    assign lfsr_next_arr[7][5] = lfsr[5] ^ lfsr[7] ^ lfsr[8] ^ lfsr[9] ^ lfsr[10] ^ lfsr[12] ^ lfsr[14] ^ lfsr[17] ^ lfsr[18] ^ lfsr[19] ^ lfsr[21] ^ lfsr[22] ^ lfsr[23] ^ lfsr[27] ^ lfsr[29] ^ lfsr[31] ^ data_i[0] ^ data_i[1] ^ data_i[3] ^ data_i[4] ^ data_i[5] ^ data_i[6] ^ data_i[7] ^ data_i[10] ^ data_i[13] ^ data_i[19] ^ data_i[20] ^ data_i[21] ^ data_i[24] ^ data_i[28] ^ data_i[29] ^ data_i[37] ^ data_i[39] ^ data_i[40] ^ data_i[41] ^ data_i[42] ^ data_i[44] ^ data_i[46] ^ data_i[49] ^ data_i[50] ^ data_i[51] ^ data_i[53] ^ data_i[54] ^ data_i[55] ^ data_i[59] ^ data_i[61] ^ data_i[63];
    assign lfsr_next_arr[7][6] = lfsr[6] ^ lfsr[8] ^ lfsr[9] ^ lfsr[10] ^ lfsr[11] ^ lfsr[13] ^ lfsr[15] ^ lfsr[18] ^ lfsr[19] ^ lfsr[20] ^ lfsr[22] ^ lfsr[23] ^ lfsr[24] ^ lfsr[28] ^ lfsr[30] ^ data_i[1] ^ data_i[2] ^ data_i[4] ^ data_i[5] ^ data_i[6] ^ data_i[7] ^ data_i[8] ^ data_i[11] ^ data_i[14] ^ data_i[20] ^ data_i[21] ^ data_i[22] ^ data_i[25] ^ data_i[29] ^ data_i[30] ^ data_i[38] ^ data_i[40] ^ data_i[41] ^ data_i[42] ^ data_i[43] ^ data_i[45] ^ data_i[47] ^ data_i[50] ^ data_i[51] ^ data_i[52] ^ data_i[54] ^ data_i[55] ^ data_i[56] ^ data_i[60] ^ data_i[62];
    assign lfsr_next_arr[7][7] = lfsr[0] ^ lfsr[2] ^ lfsr[5] ^ lfsr[7] ^ lfsr[9] ^ lfsr[10] ^ lfsr[11] ^ lfsr[13] ^ lfsr[14] ^ lfsr[15] ^ lfsr[18] ^ lfsr[19] ^ lfsr[20] ^ lfsr[22] ^ lfsr[24] ^ lfsr[25] ^ lfsr[26] ^ lfsr[28] ^ data_i[0] ^ data_i[2] ^ data_i[3] ^ data_i[5] ^ data_i[7] ^ data_i[8] ^ data_i[10] ^ data_i[15] ^ data_i[16] ^ data_i[21] ^ data_i[22] ^ data_i[23] ^ data_i[24] ^ data_i[25] ^ data_i[28] ^ data_i[29] ^ data_i[32] ^ data_i[34] ^ data_i[37] ^ data_i[39] ^ data_i[41] ^ data_i[42] ^ data_i[43] ^ data_i[45] ^ data_i[46] ^ data_i[47] ^ data_i[50] ^ data_i[51] ^ data_i[52] ^ data_i[54] ^ data_i[56] ^ data_i[57] ^ data_i[58] ^ data_i[60];
    assign lfsr_next_arr[7][8] = lfsr[0] ^ lfsr[1] ^ lfsr[2] ^ lfsr[3] ^ lfsr[5] ^ lfsr[6] ^ lfsr[8] ^ lfsr[10] ^ lfsr[11] ^ lfsr[13] ^ lfsr[14] ^ lfsr[18] ^ lfsr[19] ^ lfsr[20] ^ lfsr[22] ^ lfsr[25] ^ lfsr[27] ^ lfsr[28] ^ lfsr[31] ^ data_i[0] ^ data_i[1] ^ data_i[3] ^ data_i[4] ^ data_i[8] ^ data_i[10] ^ data_i[11] ^ data_i[12] ^ data_i[17] ^ data_i[22] ^ data_i[23] ^ data_i[28] ^ data_i[31] ^ data_i[32] ^ data_i[33] ^ data_i[34] ^ data_i[35] ^ data_i[37] ^ data_i[38] ^ data_i[40] ^ data_i[42] ^ data_i[43] ^ data_i[45] ^ data_i[46] ^ data_i[50] ^ data_i[51] ^ data_i[52] ^ data_i[54] ^ data_i[57] ^ data_i[59] ^ data_i[60] ^ data_i[63];
    assign lfsr_next_arr[7][9] = lfsr[0] ^ lfsr[1] ^ lfsr[2] ^ lfsr[3] ^ lfsr[4] ^ lfsr[6] ^ lfsr[7] ^ lfsr[9] ^ lfsr[11] ^ lfsr[12] ^ lfsr[14] ^ lfsr[15] ^ lfsr[19] ^ lfsr[20] ^ lfsr[21] ^ lfsr[23] ^ lfsr[26] ^ lfsr[28] ^ lfsr[29] ^ data_i[1] ^ data_i[2] ^ data_i[4] ^ data_i[5] ^ data_i[9] ^ data_i[11] ^ data_i[12] ^ data_i[13] ^ data_i[18] ^ data_i[23] ^ data_i[24] ^ data_i[29] ^ data_i[32] ^ data_i[33] ^ data_i[34] ^ data_i[35] ^ data_i[36] ^ data_i[38] ^ data_i[39] ^ data_i[41] ^ data_i[43] ^ data_i[44] ^ data_i[46] ^ data_i[47] ^ data_i[51] ^ data_i[52] ^ data_i[53] ^ data_i[55] ^ data_i[58] ^ data_i[60] ^ data_i[61];
    assign lfsr_next_arr[7][10] = lfsr[0] ^ lfsr[1] ^ lfsr[3] ^ lfsr[4] ^ lfsr[7] ^ lfsr[8] ^ lfsr[10] ^ lfsr[18] ^ lfsr[20] ^ lfsr[23] ^ lfsr[24] ^ lfsr[26] ^ lfsr[27] ^ lfsr[28] ^ lfsr[30] ^ lfsr[31] ^ data_i[0] ^ data_i[2] ^ data_i[3] ^ data_i[5] ^ data_i[9] ^ data_i[13] ^ data_i[14] ^ data_i[16] ^ data_i[19] ^ data_i[26] ^ data_i[28] ^ data_i[29] ^ data_i[31] ^ data_i[32] ^ data_i[33] ^ data_i[35] ^ data_i[36] ^ data_i[39] ^ data_i[40] ^ data_i[42] ^ data_i[50] ^ data_i[52] ^ data_i[55] ^ data_i[56] ^ data_i[58] ^ data_i[59] ^ data_i[60] ^ data_i[62] ^ data_i[63];
    assign lfsr_next_arr[7][11] = lfsr[1] ^ lfsr[4] ^ lfsr[8] ^ lfsr[9] ^ lfsr[11] ^ lfsr[12] ^ lfsr[13] ^ lfsr[15] ^ lfsr[16] ^ lfsr[18] ^ lfsr[19] ^ lfsr[22] ^ lfsr[23] ^ lfsr[24] ^ lfsr[25] ^ lfsr[26] ^ lfsr[27] ^ data_i[0] ^ data_i[1] ^ data_i[3] ^ data_i[4] ^ data_i[9] ^ data_i[12] ^ data_i[14] ^ data_i[15] ^ data_i[16] ^ data_i[17] ^ data_i[20] ^ data_i[24] ^ data_i[25] ^ data_i[26] ^ data_i[27] ^ data_i[28] ^ data_i[31] ^ data_i[33] ^ data_i[36] ^ data_i[40] ^ data_i[41] ^ data_i[43] ^ data_i[44] ^ data_i[45] ^ data_i[47] ^ data_i[48] ^ data_i[50] ^ data_i[51] ^ data_i[54] ^ data_i[55] ^ data_i[56] ^ data_i[57] ^ data_i[58] ^ data_i[59];
    assign lfsr_next_arr[7][12] = lfsr[9] ^ lfsr[10] ^ lfsr[14] ^ lfsr[15] ^ lfsr[17] ^ lfsr[18] ^ lfsr[19] ^ lfsr[20] ^ lfsr[21] ^ lfsr[22] ^ lfsr[24] ^ lfsr[25] ^ lfsr[27] ^ lfsr[29] ^ lfsr[31] ^ data_i[0] ^ data_i[1] ^ data_i[2] ^ data_i[4] ^ data_i[5] ^ data_i[6] ^ data_i[9] ^ data_i[12] ^ data_i[13] ^ data_i[15] ^ data_i[17] ^ data_i[18] ^ data_i[21] ^ data_i[24] ^ data_i[27] ^ data_i[30] ^ data_i[31] ^ data_i[41] ^ data_i[42] ^ data_i[46] ^ data_i[47] ^ data_i[49] ^ data_i[50] ^ data_i[51] ^ data_i[52] ^ data_i[53] ^ data_i[54] ^ data_i[56] ^ data_i[57] ^ data_i[59] ^ data_i[61] ^ data_i[63];
    assign lfsr_next_arr[7][13] = lfsr[0] ^ lfsr[10] ^ lfsr[11] ^ lfsr[15] ^ lfsr[16] ^ lfsr[18] ^ lfsr[19] ^ lfsr[20] ^ lfsr[21] ^ lfsr[22] ^ lfsr[23] ^ lfsr[25] ^ lfsr[26] ^ lfsr[28] ^ lfsr[30] ^ data_i[1] ^ data_i[2] ^ data_i[3] ^ data_i[5] ^ data_i[6] ^ data_i[7] ^ data_i[10] ^ data_i[13] ^ data_i[14] ^ data_i[16] ^ data_i[18] ^ data_i[19] ^ data_i[22] ^ data_i[25] ^ data_i[28] ^ data_i[31] ^ data_i[32] ^ data_i[42] ^ data_i[43] ^ data_i[47] ^ data_i[48] ^ data_i[50] ^ data_i[51] ^ data_i[52] ^ data_i[53] ^ data_i[54] ^ data_i[55] ^ data_i[57] ^ data_i[58] ^ data_i[60] ^ data_i[62];
    assign lfsr_next_arr[7][14] = lfsr[0] ^ lfsr[1] ^ lfsr[11] ^ lfsr[12] ^ lfsr[16] ^ lfsr[17] ^ lfsr[19] ^ lfsr[20] ^ lfsr[21] ^ lfsr[22] ^ lfsr[23] ^ lfsr[24] ^ lfsr[26] ^ lfsr[27] ^ lfsr[29] ^ lfsr[31] ^ data_i[2] ^ data_i[3] ^ data_i[4] ^ data_i[6] ^ data_i[7] ^ data_i[8] ^ data_i[11] ^ data_i[14] ^ data_i[15] ^ data_i[17] ^ data_i[19] ^ data_i[20] ^ data_i[23] ^ data_i[26] ^ data_i[29] ^ data_i[32] ^ data_i[33] ^ data_i[43] ^ data_i[44] ^ data_i[48] ^ data_i[49] ^ data_i[51] ^ data_i[52] ^ data_i[53] ^ data_i[54] ^ data_i[55] ^ data_i[56] ^ data_i[58] ^ data_i[59] ^ data_i[61] ^ data_i[63];
    assign lfsr_next_arr[7][15] = lfsr[1] ^ lfsr[2] ^ lfsr[12] ^ lfsr[13] ^ lfsr[17] ^ lfsr[18] ^ lfsr[20] ^ lfsr[21] ^ lfsr[22] ^ lfsr[23] ^ lfsr[24] ^ lfsr[25] ^ lfsr[27] ^ lfsr[28] ^ lfsr[30] ^ data_i[3] ^ data_i[4] ^ data_i[5] ^ data_i[7] ^ data_i[8] ^ data_i[9] ^ data_i[12] ^ data_i[15] ^ data_i[16] ^ data_i[18] ^ data_i[20] ^ data_i[21] ^ data_i[24] ^ data_i[27] ^ data_i[30] ^ data_i[33] ^ data_i[34] ^ data_i[44] ^ data_i[45] ^ data_i[49] ^ data_i[50] ^ data_i[52] ^ data_i[53] ^ data_i[54] ^ data_i[55] ^ data_i[56] ^ data_i[57] ^ data_i[59] ^ data_i[60] ^ data_i[62];
    assign lfsr_next_arr[7][16] = lfsr[0] ^ lfsr[3] ^ lfsr[5] ^ lfsr[12] ^ lfsr[14] ^ lfsr[15] ^ lfsr[16] ^ lfsr[19] ^ lfsr[24] ^ lfsr[25] ^ data_i[0] ^ data_i[4] ^ data_i[5] ^ data_i[8] ^ data_i[12] ^ data_i[13] ^ data_i[17] ^ data_i[19] ^ data_i[21] ^ data_i[22] ^ data_i[24] ^ data_i[26] ^ data_i[29] ^ data_i[30] ^ data_i[32] ^ data_i[35] ^ data_i[37] ^ data_i[44] ^ data_i[46] ^ data_i[47] ^ data_i[48] ^ data_i[51] ^ data_i[56] ^ data_i[57];
    assign lfsr_next_arr[7][17] = lfsr[1] ^ lfsr[4] ^ lfsr[6] ^ lfsr[13] ^ lfsr[15] ^ lfsr[16] ^ lfsr[17] ^ lfsr[20] ^ lfsr[25] ^ lfsr[26] ^ data_i[1] ^ data_i[5] ^ data_i[6] ^ data_i[9] ^ data_i[13] ^ data_i[14] ^ data_i[18] ^ data_i[20] ^ data_i[22] ^ data_i[23] ^ data_i[25] ^ data_i[27] ^ data_i[30] ^ data_i[31] ^ data_i[33] ^ data_i[36] ^ data_i[38] ^ data_i[45] ^ data_i[47] ^ data_i[48] ^ data_i[49] ^ data_i[52] ^ data_i[57] ^ data_i[58];
    assign lfsr_next_arr[7][18] = lfsr[0] ^ lfsr[2] ^ lfsr[5] ^ lfsr[7] ^ lfsr[14] ^ lfsr[16] ^ lfsr[17] ^ lfsr[18] ^ lfsr[21] ^ lfsr[26] ^ lfsr[27] ^ data_i[2] ^ data_i[6] ^ data_i[7] ^ data_i[10] ^ data_i[14] ^ data_i[15] ^ data_i[19] ^ data_i[21] ^ data_i[23] ^ data_i[24] ^ data_i[26] ^ data_i[28] ^ data_i[31] ^ data_i[32] ^ data_i[34] ^ data_i[37] ^ data_i[39] ^ data_i[46] ^ data_i[48] ^ data_i[49] ^ data_i[50] ^ data_i[53] ^ data_i[58] ^ data_i[59];
    assign lfsr_next_arr[7][19] = lfsr[0] ^ lfsr[1] ^ lfsr[3] ^ lfsr[6] ^ lfsr[8] ^ lfsr[15] ^ lfsr[17] ^ lfsr[18] ^ lfsr[19] ^ lfsr[22] ^ lfsr[27] ^ lfsr[28] ^ data_i[3] ^ data_i[7] ^ data_i[8] ^ data_i[11] ^ data_i[15] ^ data_i[16] ^ data_i[20] ^ data_i[22] ^ data_i[24] ^ data_i[25] ^ data_i[27] ^ data_i[29] ^ data_i[32] ^ data_i[33] ^ data_i[35] ^ data_i[38] ^ data_i[40] ^ data_i[47] ^ data_i[49] ^ data_i[50] ^ data_i[51] ^ data_i[54] ^ data_i[59] ^ data_i[60];
    assign lfsr_next_arr[7][20] = lfsr[1] ^ lfsr[2] ^ lfsr[4] ^ lfsr[7] ^ lfsr[9] ^ lfsr[16] ^ lfsr[18] ^ lfsr[19] ^ lfsr[20] ^ lfsr[23] ^ lfsr[28] ^ lfsr[29] ^ data_i[4] ^ data_i[8] ^ data_i[9] ^ data_i[12] ^ data_i[16] ^ data_i[17] ^ data_i[21] ^ data_i[23] ^ data_i[25] ^ data_i[26] ^ data_i[28] ^ data_i[30] ^ data_i[33] ^ data_i[34] ^ data_i[36] ^ data_i[39] ^ data_i[41] ^ data_i[48] ^ data_i[50] ^ data_i[51] ^ data_i[52] ^ data_i[55] ^ data_i[60] ^ data_i[61];
    assign lfsr_next_arr[7][21] = lfsr[2] ^ lfsr[3] ^ lfsr[5] ^ lfsr[8] ^ lfsr[10] ^ lfsr[17] ^ lfsr[19] ^ lfsr[20] ^ lfsr[21] ^ lfsr[24] ^ lfsr[29] ^ lfsr[30] ^ data_i[5] ^ data_i[9] ^ data_i[10] ^ data_i[13] ^ data_i[17] ^ data_i[18] ^ data_i[22] ^ data_i[24] ^ data_i[26] ^ data_i[27] ^ data_i[29] ^ data_i[31] ^ data_i[34] ^ data_i[35] ^ data_i[37] ^ data_i[40] ^ data_i[42] ^ data_i[49] ^ data_i[51] ^ data_i[52] ^ data_i[53] ^ data_i[56] ^ data_i[61] ^ data_i[62];
    assign lfsr_next_arr[7][22] = lfsr[2] ^ lfsr[3] ^ lfsr[4] ^ lfsr[5] ^ lfsr[6] ^ lfsr[9] ^ lfsr[11] ^ lfsr[12] ^ lfsr[13] ^ lfsr[15] ^ lfsr[16] ^ lfsr[20] ^ lfsr[23] ^ lfsr[25] ^ lfsr[26] ^ lfsr[28] ^ lfsr[29] ^ lfsr[30] ^ data_i[0] ^ data_i[9] ^ data_i[11] ^ data_i[12] ^ data_i[14] ^ data_i[16] ^ data_i[18] ^ data_i[19] ^ data_i[23] ^ data_i[24] ^ data_i[26] ^ data_i[27] ^ data_i[29] ^ data_i[31] ^ data_i[34] ^ data_i[35] ^ data_i[36] ^ data_i[37] ^ data_i[38] ^ data_i[41] ^ data_i[43] ^ data_i[44] ^ data_i[45] ^ data_i[47] ^ data_i[48] ^ data_i[52] ^ data_i[55] ^ data_i[57] ^ data_i[58] ^ data_i[60] ^ data_i[61] ^ data_i[62];
    assign lfsr_next_arr[7][23] = lfsr[2] ^ lfsr[3] ^ lfsr[4] ^ lfsr[6] ^ lfsr[7] ^ lfsr[10] ^ lfsr[14] ^ lfsr[15] ^ lfsr[17] ^ lfsr[18] ^ lfsr[22] ^ lfsr[23] ^ lfsr[24] ^ lfsr[27] ^ lfsr[28] ^ lfsr[30] ^ data_i[0] ^ data_i[1] ^ data_i[6] ^ data_i[9] ^ data_i[13] ^ data_i[15] ^ data_i[16] ^ data_i[17] ^ data_i[19] ^ data_i[20] ^ data_i[26] ^ data_i[27] ^ data_i[29] ^ data_i[31] ^ data_i[34] ^ data_i[35] ^ data_i[36] ^ data_i[38] ^ data_i[39] ^ data_i[42] ^ data_i[46] ^ data_i[47] ^ data_i[49] ^ data_i[50] ^ data_i[54] ^ data_i[55] ^ data_i[56] ^ data_i[59] ^ data_i[60] ^ data_i[62];
    assign lfsr_next_arr[7][24] = lfsr[0] ^ lfsr[3] ^ lfsr[4] ^ lfsr[5] ^ lfsr[7] ^ lfsr[8] ^ lfsr[11] ^ lfsr[15] ^ lfsr[16] ^ lfsr[18] ^ lfsr[19] ^ lfsr[23] ^ lfsr[24] ^ lfsr[25] ^ lfsr[28] ^ lfsr[29] ^ lfsr[31] ^ data_i[1] ^ data_i[2] ^ data_i[7] ^ data_i[10] ^ data_i[14] ^ data_i[16] ^ data_i[17] ^ data_i[18] ^ data_i[20] ^ data_i[21] ^ data_i[27] ^ data_i[28] ^ data_i[30] ^ data_i[32] ^ data_i[35] ^ data_i[36] ^ data_i[37] ^ data_i[39] ^ data_i[40] ^ data_i[43] ^ data_i[47] ^ data_i[48] ^ data_i[50] ^ data_i[51] ^ data_i[55] ^ data_i[56] ^ data_i[57] ^ data_i[60] ^ data_i[61] ^ data_i[63];
    assign lfsr_next_arr[7][25] = lfsr[1] ^ lfsr[4] ^ lfsr[5] ^ lfsr[6] ^ lfsr[8] ^ lfsr[9] ^ lfsr[12] ^ lfsr[16] ^ lfsr[17] ^ lfsr[19] ^ lfsr[20] ^ lfsr[24] ^ lfsr[25] ^ lfsr[26] ^ lfsr[29] ^ lfsr[30] ^ data_i[2] ^ data_i[3] ^ data_i[8] ^ data_i[11] ^ data_i[15] ^ data_i[17] ^ data_i[18] ^ data_i[19] ^ data_i[21] ^ data_i[22] ^ data_i[28] ^ data_i[29] ^ data_i[31] ^ data_i[33] ^ data_i[36] ^ data_i[37] ^ data_i[38] ^ data_i[40] ^ data_i[41] ^ data_i[44] ^ data_i[48] ^ data_i[49] ^ data_i[51] ^ data_i[52] ^ data_i[56] ^ data_i[57] ^ data_i[58] ^ data_i[61] ^ data_i[62];
    assign lfsr_next_arr[7][26] = lfsr[6] ^ lfsr[7] ^ lfsr[9] ^ lfsr[10] ^ lfsr[12] ^ lfsr[15] ^ lfsr[16] ^ lfsr[17] ^ lfsr[20] ^ lfsr[22] ^ lfsr[23] ^ lfsr[25] ^ lfsr[27] ^ lfsr[28] ^ lfsr[29] ^ lfsr[30] ^ data_i[0] ^ data_i[3] ^ data_i[4] ^ data_i[6] ^ data_i[10] ^ data_i[18] ^ data_i[19] ^ data_i[20] ^ data_i[22] ^ data_i[23] ^ data_i[24] ^ data_i[25] ^ data_i[26] ^ data_i[28] ^ data_i[31] ^ data_i[38] ^ data_i[39] ^ data_i[41] ^ data_i[42] ^ data_i[44] ^ data_i[47] ^ data_i[48] ^ data_i[49] ^ data_i[52] ^ data_i[54] ^ data_i[55] ^ data_i[57] ^ data_i[59] ^ data_i[60] ^ data_i[61] ^ data_i[62];
    assign lfsr_next_arr[7][27] = lfsr[0] ^ lfsr[7] ^ lfsr[8] ^ lfsr[10] ^ lfsr[11] ^ lfsr[13] ^ lfsr[16] ^ lfsr[17] ^ lfsr[18] ^ lfsr[21] ^ lfsr[23] ^ lfsr[24] ^ lfsr[26] ^ lfsr[28] ^ lfsr[29] ^ lfsr[30] ^ lfsr[31] ^ data_i[1] ^ data_i[4] ^ data_i[5] ^ data_i[7] ^ data_i[11] ^ data_i[19] ^ data_i[20] ^ data_i[21] ^ data_i[23] ^ data_i[24] ^ data_i[25] ^ data_i[26] ^ data_i[27] ^ data_i[29] ^ data_i[32] ^ data_i[39] ^ data_i[40] ^ data_i[42] ^ data_i[43] ^ data_i[45] ^ data_i[48] ^ data_i[49] ^ data_i[50] ^ data_i[53] ^ data_i[55] ^ data_i[56] ^ data_i[58] ^ data_i[60] ^ data_i[61] ^ data_i[62] ^ data_i[63];
    assign lfsr_next_arr[7][28] = lfsr[1] ^ lfsr[8] ^ lfsr[9] ^ lfsr[11] ^ lfsr[12] ^ lfsr[14] ^ lfsr[17] ^ lfsr[18] ^ lfsr[19] ^ lfsr[22] ^ lfsr[24] ^ lfsr[25] ^ lfsr[27] ^ lfsr[29] ^ lfsr[30] ^ lfsr[31] ^ data_i[2] ^ data_i[5] ^ data_i[6] ^ data_i[8] ^ data_i[12] ^ data_i[20] ^ data_i[21] ^ data_i[22] ^ data_i[24] ^ data_i[25] ^ data_i[26] ^ data_i[27] ^ data_i[28] ^ data_i[30] ^ data_i[33] ^ data_i[40] ^ data_i[41] ^ data_i[43] ^ data_i[44] ^ data_i[46] ^ data_i[49] ^ data_i[50] ^ data_i[51] ^ data_i[54] ^ data_i[56] ^ data_i[57] ^ data_i[59] ^ data_i[61] ^ data_i[62] ^ data_i[63];
    assign lfsr_next_arr[7][29] = lfsr[2] ^ lfsr[9] ^ lfsr[10] ^ lfsr[12] ^ lfsr[13] ^ lfsr[15] ^ lfsr[18] ^ lfsr[19] ^ lfsr[20] ^ lfsr[23] ^ lfsr[25] ^ lfsr[26] ^ lfsr[28] ^ lfsr[30] ^ lfsr[31] ^ data_i[3] ^ data_i[6] ^ data_i[7] ^ data_i[9] ^ data_i[13] ^ data_i[21] ^ data_i[22] ^ data_i[23] ^ data_i[25] ^ data_i[26] ^ data_i[27] ^ data_i[28] ^ data_i[29] ^ data_i[31] ^ data_i[34] ^ data_i[41] ^ data_i[42] ^ data_i[44] ^ data_i[45] ^ data_i[47] ^ data_i[50] ^ data_i[51] ^ data_i[52] ^ data_i[55] ^ data_i[57] ^ data_i[58] ^ data_i[60] ^ data_i[62] ^ data_i[63];
    assign lfsr_next_arr[7][30] = lfsr[0] ^ lfsr[3] ^ lfsr[10] ^ lfsr[11] ^ lfsr[13] ^ lfsr[14] ^ lfsr[16] ^ lfsr[19] ^ lfsr[20] ^ lfsr[21] ^ lfsr[24] ^ lfsr[26] ^ lfsr[27] ^ lfsr[29] ^ lfsr[31] ^ data_i[4] ^ data_i[7] ^ data_i[8] ^ data_i[10] ^ data_i[14] ^ data_i[22] ^ data_i[23] ^ data_i[24] ^ data_i[26] ^ data_i[27] ^ data_i[28] ^ data_i[29] ^ data_i[30] ^ data_i[32] ^ data_i[35] ^ data_i[42] ^ data_i[43] ^ data_i[45] ^ data_i[46] ^ data_i[48] ^ data_i[51] ^ data_i[52] ^ data_i[53] ^ data_i[56] ^ data_i[58] ^ data_i[59] ^ data_i[61] ^ data_i[63];
    assign lfsr_next_arr[7][31] = lfsr[1] ^ lfsr[4] ^ lfsr[11] ^ lfsr[12] ^ lfsr[14] ^ lfsr[15] ^ lfsr[17] ^ lfsr[20] ^ lfsr[21] ^ lfsr[22] ^ lfsr[25] ^ lfsr[27] ^ lfsr[28] ^ lfsr[30] ^ data_i[5] ^ data_i[8] ^ data_i[9] ^ data_i[11] ^ data_i[15] ^ data_i[23] ^ data_i[24] ^ data_i[25] ^ data_i[27] ^ data_i[28] ^ data_i[29] ^ data_i[30] ^ data_i[31] ^ data_i[33] ^ data_i[36] ^ data_i[43] ^ data_i[44] ^ data_i[46] ^ data_i[47] ^ data_i[49] ^ data_i[52] ^ data_i[53] ^ data_i[54] ^ data_i[57] ^ data_i[59] ^ data_i[60] ^ data_i[62];
end

/* select next lfst based on number of valid bytes */
always_comb begin
	for(int i=0; i<KEEP_W; i++) begin : crc_lfsr_loop
		/* verilator lint_off WIDTHEXPAND */
		if( (i+1) == len_i )lfsr_next = lfsr_next_arr[i];
		/* verilator lint_on WIDTHEXPAND */
	end
end

  always @(posedge clk) begin
    if ( valid_i )  begin
      lfsr_q <= lfsr_next;
    end
  end // always
endmodule // crc
