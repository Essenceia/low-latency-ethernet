module tcp_client(
);

endmodule
