//-----------------------------------------------------------------------------
// Copyright (C) 2009 OutputLogic.com
// This source file may be used and distributed without restriction
// provided that this copyright statement is not removed from the file
// and that any derivative work contains the original copyright notice
// and the associated disclaimer.
//
// THIS SOURCE FILE IS PROVIDED "AS IS" AND WITHOUT ANY EXPRESS
// OR IMPLIED WARRANTIES, INCLUDING, WITHOUT LIMITATION, THE IMPLIED
// WARRANTIES OF MERCHANTIBILITY AND FITNESS FOR A PARTICULAR PURPOSE.
//-----------------------------------------------------------------------------
// CRC module for data[31:0] ,   crc[31:0]=1+x^1+x^2+x^4+x^5+x^7+x^8+x^10+x^11+x^12+x^16+x^22+x^23+x^26+x^32;
//-----------------------------------------------------------------------------
module crc #(
	parameter DATA_W = 32,
	parameter CRC_W = 32
)
(
  input               clk,
  input               valid_i,
  input               start_i,
  input  [DATA_W-1:0] data_i,
  output [CRC_W-1:0]  crc_o
);

  reg   [CRC_W-1:0] lfsr_q;
  logic [CRC_W-1:0] lfsr_next;
  logic [CRC_W-1:0] lfsr;

  assign crc_o = lfsr_q;
  assign lfsr = start_i ? {CRC_W{1'b1}} : lfsr_q;

if(DATA_W == 16) begin
  assign  lfsr_next[0] = lfsr[16] ^ lfsr[22] ^ lfsr[25] ^ lfsr[26] ^ lfsr[28] ^ data_i[0] ^ data_i[6] ^ data_i[9] ^ data_i[10] ^ data_i[12];
  assign  lfsr_next[1] = lfsr[16] ^ lfsr[17] ^ lfsr[22] ^ lfsr[23] ^ lfsr[25] ^ lfsr[27] ^ lfsr[28] ^ lfsr[29] ^ data_i[0] ^ data_i[1] ^ data_i[6] ^ data_i[7] ^ data_i[9] ^ data_i[11] ^ data_i[12] ^ data_i[13];
  assign  lfsr_next[2] = lfsr[16] ^ lfsr[17] ^ lfsr[18] ^ lfsr[22] ^ lfsr[23] ^ lfsr[24] ^ lfsr[25] ^ lfsr[29] ^ lfsr[30] ^ data_i[0] ^ data_i[1] ^ data_i[2] ^ data_i[6] ^ data_i[7] ^ data_i[8] ^ data_i[9] ^ data_i[13] ^ data_i[14];
  assign  lfsr_next[3] = lfsr[17] ^ lfsr[18] ^ lfsr[19] ^ lfsr[23] ^ lfsr[24] ^ lfsr[25] ^ lfsr[26] ^ lfsr[30] ^ lfsr[31] ^ data_i[1] ^ data_i[2] ^ data_i[3] ^ data_i[7] ^ data_i[8] ^ data_i[9] ^ data_i[10] ^ data_i[14] ^ data_i[15];
  assign  lfsr_next[4] = lfsr[16] ^ lfsr[18] ^ lfsr[19] ^ lfsr[20] ^ lfsr[22] ^ lfsr[24] ^ lfsr[27] ^ lfsr[28] ^ lfsr[31] ^ data_i[0] ^ data_i[2] ^ data_i[3] ^ data_i[4] ^ data_i[6] ^ data_i[8] ^ data_i[11] ^ data_i[12] ^ data_i[15];
  assign  lfsr_next[5] = lfsr[16] ^ lfsr[17] ^ lfsr[19] ^ lfsr[20] ^ lfsr[21] ^ lfsr[22] ^ lfsr[23] ^ lfsr[26] ^ lfsr[29] ^ data_i[0] ^ data_i[1] ^ data_i[3] ^ data_i[4] ^ data_i[5] ^ data_i[6] ^ data_i[7] ^ data_i[10] ^ data_i[13];
  assign  lfsr_next[6] = lfsr[17] ^ lfsr[18] ^ lfsr[20] ^ lfsr[21] ^ lfsr[22] ^ lfsr[23] ^ lfsr[24] ^ lfsr[27] ^ lfsr[30] ^ data_i[1] ^ data_i[2] ^ data_i[4] ^ data_i[5] ^ data_i[6] ^ data_i[7] ^ data_i[8] ^ data_i[11] ^ data_i[14];
  assign  lfsr_next[7] = lfsr[16] ^ lfsr[18] ^ lfsr[19] ^ lfsr[21] ^ lfsr[23] ^ lfsr[24] ^ lfsr[26] ^ lfsr[31] ^ data_i[0] ^ data_i[2] ^ data_i[3] ^ data_i[5] ^ data_i[7] ^ data_i[8] ^ data_i[10] ^ data_i[15];
  assign  lfsr_next[8] = lfsr[16] ^ lfsr[17] ^ lfsr[19] ^ lfsr[20] ^ lfsr[24] ^ lfsr[26] ^ lfsr[27] ^ lfsr[28] ^ data_i[0] ^ data_i[1] ^ data_i[3] ^ data_i[4] ^ data_i[8] ^ data_i[10] ^ data_i[11] ^ data_i[12];
  assign  lfsr_next[9] = lfsr[17] ^ lfsr[18] ^ lfsr[20] ^ lfsr[21] ^ lfsr[25] ^ lfsr[27] ^ lfsr[28] ^ lfsr[29] ^ data_i[1] ^ data_i[2] ^ data_i[4] ^ data_i[5] ^ data_i[9] ^ data_i[11] ^ data_i[12] ^ data_i[13];
  assign  lfsr_next[10] = lfsr[16] ^ lfsr[18] ^ lfsr[19] ^ lfsr[21] ^ lfsr[25] ^ lfsr[29] ^ lfsr[30] ^ data_i[0] ^ data_i[2] ^ data_i[3] ^ data_i[5] ^ data_i[9] ^ data_i[13] ^ data_i[14];
  assign  lfsr_next[11] = lfsr[16] ^ lfsr[17] ^ lfsr[19] ^ lfsr[20] ^ lfsr[25] ^ lfsr[28] ^ lfsr[30] ^ lfsr[31] ^ data_i[0] ^ data_i[1] ^ data_i[3] ^ data_i[4] ^ data_i[9] ^ data_i[12] ^ data_i[14] ^ data_i[15];
  assign  lfsr_next[12] = lfsr[16] ^ lfsr[17] ^ lfsr[18] ^ lfsr[20] ^ lfsr[21] ^ lfsr[22] ^ lfsr[25] ^ lfsr[28] ^ lfsr[29] ^ lfsr[31] ^ data_i[0] ^ data_i[1] ^ data_i[2] ^ data_i[4] ^ data_i[5] ^ data_i[6] ^ data_i[9] ^ data_i[12] ^ data_i[13] ^ data_i[15];
  assign  lfsr_next[13] = lfsr[17] ^ lfsr[18] ^ lfsr[19] ^ lfsr[21] ^ lfsr[22] ^ lfsr[23] ^ lfsr[26] ^ lfsr[29] ^ lfsr[30] ^ data_i[1] ^ data_i[2] ^ data_i[3] ^ data_i[5] ^ data_i[6] ^ data_i[7] ^ data_i[10] ^ data_i[13] ^ data_i[14];
  assign  lfsr_next[14] = lfsr[18] ^ lfsr[19] ^ lfsr[20] ^ lfsr[22] ^ lfsr[23] ^ lfsr[24] ^ lfsr[27] ^ lfsr[30] ^ lfsr[31] ^ data_i[2] ^ data_i[3] ^ data_i[4] ^ data_i[6] ^ data_i[7] ^ data_i[8] ^ data_i[11] ^ data_i[14] ^ data_i[15];
  assign  lfsr_next[15] = lfsr[19] ^ lfsr[20] ^ lfsr[21] ^ lfsr[23] ^ lfsr[24] ^ lfsr[25] ^ lfsr[28] ^ lfsr[31] ^ data_i[3] ^ data_i[4] ^ data_i[5] ^ data_i[7] ^ data_i[8] ^ data_i[9] ^ data_i[12] ^ data_i[15];
  assign  lfsr_next[16] = lfsr[0] ^ lfsr[16] ^ lfsr[20] ^ lfsr[21] ^ lfsr[24] ^ lfsr[28] ^ lfsr[29] ^ data_i[0] ^ data_i[4] ^ data_i[5] ^ data_i[8] ^ data_i[12] ^ data_i[13];
  assign  lfsr_next[17] = lfsr[1] ^ lfsr[17] ^ lfsr[21] ^ lfsr[22] ^ lfsr[25] ^ lfsr[29] ^ lfsr[30] ^ data_i[1] ^ data_i[5] ^ data_i[6] ^ data_i[9] ^ data_i[13] ^ data_i[14];
  assign  lfsr_next[18] = lfsr[2] ^ lfsr[18] ^ lfsr[22] ^ lfsr[23] ^ lfsr[26] ^ lfsr[30] ^ lfsr[31] ^ data_i[2] ^ data_i[6] ^ data_i[7] ^ data_i[10] ^ data_i[14] ^ data_i[15];
  assign  lfsr_next[19] = lfsr[3] ^ lfsr[19] ^ lfsr[23] ^ lfsr[24] ^ lfsr[27] ^ lfsr[31] ^ data_i[3] ^ data_i[7] ^ data_i[8] ^ data_i[11] ^ data_i[15];
  assign  lfsr_next[20] = lfsr[4] ^ lfsr[20] ^ lfsr[24] ^ lfsr[25] ^ lfsr[28] ^ data_i[4] ^ data_i[8] ^ data_i[9] ^ data_i[12];
  assign  lfsr_next[21] = lfsr[5] ^ lfsr[21] ^ lfsr[25] ^ lfsr[26] ^ lfsr[29] ^ data_i[5] ^ data_i[9] ^ data_i[10] ^ data_i[13];
  assign  lfsr_next[22] = lfsr[6] ^ lfsr[16] ^ lfsr[25] ^ lfsr[27] ^ lfsr[28] ^ lfsr[30] ^ data_i[0] ^ data_i[9] ^ data_i[11] ^ data_i[12] ^ data_i[14];
  assign  lfsr_next[23] = lfsr[7] ^ lfsr[16] ^ lfsr[17] ^ lfsr[22] ^ lfsr[25] ^ lfsr[29] ^ lfsr[31] ^ data_i[0] ^ data_i[1] ^ data_i[6] ^ data_i[9] ^ data_i[13] ^ data_i[15];
  assign  lfsr_next[24] = lfsr[8] ^ lfsr[17] ^ lfsr[18] ^ lfsr[23] ^ lfsr[26] ^ lfsr[30] ^ data_i[1] ^ data_i[2] ^ data_i[7] ^ data_i[10] ^ data_i[14];
  assign  lfsr_next[25] = lfsr[9] ^ lfsr[18] ^ lfsr[19] ^ lfsr[24] ^ lfsr[27] ^ lfsr[31] ^ data_i[2] ^ data_i[3] ^ data_i[8] ^ data_i[11] ^ data_i[15];
  assign  lfsr_next[26] = lfsr[10] ^ lfsr[16] ^ lfsr[19] ^ lfsr[20] ^ lfsr[22] ^ lfsr[26] ^ data_i[0] ^ data_i[3] ^ data_i[4] ^ data_i[6] ^ data_i[10];
  assign  lfsr_next[27] = lfsr[11] ^ lfsr[17] ^ lfsr[20] ^ lfsr[21] ^ lfsr[23] ^ lfsr[27] ^ data_i[1] ^ data_i[4] ^ data_i[5] ^ data_i[7] ^ data_i[11];
  assign  lfsr_next[28] = lfsr[12] ^ lfsr[18] ^ lfsr[21] ^ lfsr[22] ^ lfsr[24] ^ lfsr[28] ^ data_i[2] ^ data_i[5] ^ data_i[6] ^ data_i[8] ^ data_i[12];
  assign  lfsr_next[29] = lfsr[13] ^ lfsr[19] ^ lfsr[22] ^ lfsr[23] ^ lfsr[25] ^ lfsr[29] ^ data_i[3] ^ data_i[6] ^ data_i[7] ^ data_i[9] ^ data_i[13];
  assign  lfsr_next[30] = lfsr[14] ^ lfsr[20] ^ lfsr[23] ^ lfsr[24] ^ lfsr[26] ^ lfsr[30] ^ data_i[4] ^ data_i[7] ^ data_i[8] ^ data_i[10] ^ data_i[14];
  assign  lfsr_next[31] = lfsr[15] ^ lfsr[21] ^ lfsr[24] ^ lfsr[25] ^ lfsr[27] ^ lfsr[31] ^ data_i[5] ^ data_i[8] ^ data_i[9] ^ data_i[11] ^ data_i[15];
end else if(DATA_W == 32) begin
   assign lfsr_next[0] = lfsr[0] ^ lfsr[6] ^ lfsr[9] ^ lfsr[10] ^ lfsr[12] ^ lfsr[16] ^ lfsr[24] ^ lfsr[25] ^ lfsr[26] ^ lfsr[28] ^ lfsr[29] ^ lfsr[30] ^ lfsr[31] ^ data_i[0] ^ data_i[6] ^ data_i[9] ^ data_i[10] ^ data_i[12] ^ data_i[16] ^ data_i[24] ^ data_i[25] ^ data_i[26] ^ data_i[28] ^ data_i[29] ^ data_i[30] ^ data_i[31];
   assign lfsr_next[1] = lfsr[0] ^ lfsr[1] ^ lfsr[6] ^ lfsr[7] ^ lfsr[9] ^ lfsr[11] ^ lfsr[12] ^ lfsr[13] ^ lfsr[16] ^ lfsr[17] ^ lfsr[24] ^ lfsr[27] ^ lfsr[28] ^ data_i[0] ^ data_i[1] ^ data_i[6] ^ data_i[7] ^ data_i[9] ^ data_i[11] ^ data_i[12] ^ data_i[13] ^ data_i[16] ^ data_i[17] ^ data_i[24] ^ data_i[27] ^ data_i[28];
   assign lfsr_next[2] = lfsr[0] ^ lfsr[1] ^ lfsr[2] ^ lfsr[6] ^ lfsr[7] ^ lfsr[8] ^ lfsr[9] ^ lfsr[13] ^ lfsr[14] ^ lfsr[16] ^ lfsr[17] ^ lfsr[18] ^ lfsr[24] ^ lfsr[26] ^ lfsr[30] ^ lfsr[31] ^ data_i[0] ^ data_i[1] ^ data_i[2] ^ data_i[6] ^ data_i[7] ^ data_i[8] ^ data_i[9] ^ data_i[13] ^ data_i[14] ^ data_i[16] ^ data_i[17] ^ data_i[18] ^ data_i[24] ^ data_i[26] ^ data_i[30] ^ data_i[31];
   assign lfsr_next[3] = lfsr[1] ^ lfsr[2] ^ lfsr[3] ^ lfsr[7] ^ lfsr[8] ^ lfsr[9] ^ lfsr[10] ^ lfsr[14] ^ lfsr[15] ^ lfsr[17] ^ lfsr[18] ^ lfsr[19] ^ lfsr[25] ^ lfsr[27] ^ lfsr[31] ^ data_i[1] ^ data_i[2] ^ data_i[3] ^ data_i[7] ^ data_i[8] ^ data_i[9] ^ data_i[10] ^ data_i[14] ^ data_i[15] ^ data_i[17] ^ data_i[18] ^ data_i[19] ^ data_i[25] ^ data_i[27] ^ data_i[31];
   assign lfsr_next[4] = lfsr[0] ^ lfsr[2] ^ lfsr[3] ^ lfsr[4] ^ lfsr[6] ^ lfsr[8] ^ lfsr[11] ^ lfsr[12] ^ lfsr[15] ^ lfsr[18] ^ lfsr[19] ^ lfsr[20] ^ lfsr[24] ^ lfsr[25] ^ lfsr[29] ^ lfsr[30] ^ lfsr[31] ^ data_i[0] ^ data_i[2] ^ data_i[3] ^ data_i[4] ^ data_i[6] ^ data_i[8] ^ data_i[11] ^ data_i[12] ^ data_i[15] ^ data_i[18] ^ data_i[19] ^ data_i[20] ^ data_i[24] ^ data_i[25] ^ data_i[29] ^ data_i[30] ^ data_i[31];
   assign lfsr_next[5] = lfsr[0] ^ lfsr[1] ^ lfsr[3] ^ lfsr[4] ^ lfsr[5] ^ lfsr[6] ^ lfsr[7] ^ lfsr[10] ^ lfsr[13] ^ lfsr[19] ^ lfsr[20] ^ lfsr[21] ^ lfsr[24] ^ lfsr[28] ^ lfsr[29] ^ data_i[0] ^ data_i[1] ^ data_i[3] ^ data_i[4] ^ data_i[5] ^ data_i[6] ^ data_i[7] ^ data_i[10] ^ data_i[13] ^ data_i[19] ^ data_i[20] ^ data_i[21] ^ data_i[24] ^ data_i[28] ^ data_i[29];
   assign lfsr_next[6] = lfsr[1] ^ lfsr[2] ^ lfsr[4] ^ lfsr[5] ^ lfsr[6] ^ lfsr[7] ^ lfsr[8] ^ lfsr[11] ^ lfsr[14] ^ lfsr[20] ^ lfsr[21] ^ lfsr[22] ^ lfsr[25] ^ lfsr[29] ^ lfsr[30] ^ data_i[1] ^ data_i[2] ^ data_i[4] ^ data_i[5] ^ data_i[6] ^ data_i[7] ^ data_i[8] ^ data_i[11] ^ data_i[14] ^ data_i[20] ^ data_i[21] ^ data_i[22] ^ data_i[25] ^ data_i[29] ^ data_i[30];
   assign lfsr_next[7] = lfsr[0] ^ lfsr[2] ^ lfsr[3] ^ lfsr[5] ^ lfsr[7] ^ lfsr[8] ^ lfsr[10] ^ lfsr[15] ^ lfsr[16] ^ lfsr[21] ^ lfsr[22] ^ lfsr[23] ^ lfsr[24] ^ lfsr[25] ^ lfsr[28] ^ lfsr[29] ^ data_i[0] ^ data_i[2] ^ data_i[3] ^ data_i[5] ^ data_i[7] ^ data_i[8] ^ data_i[10] ^ data_i[15] ^ data_i[16] ^ data_i[21] ^ data_i[22] ^ data_i[23] ^ data_i[24] ^ data_i[25] ^ data_i[28] ^ data_i[29];
   assign lfsr_next[8] = lfsr[0] ^ lfsr[1] ^ lfsr[3] ^ lfsr[4] ^ lfsr[8] ^ lfsr[10] ^ lfsr[11] ^ lfsr[12] ^ lfsr[17] ^ lfsr[22] ^ lfsr[23] ^ lfsr[28] ^ lfsr[31] ^ data_i[0] ^ data_i[1] ^ data_i[3] ^ data_i[4] ^ data_i[8] ^ data_i[10] ^ data_i[11] ^ data_i[12] ^ data_i[17] ^ data_i[22] ^ data_i[23] ^ data_i[28] ^ data_i[31];
   assign lfsr_next[9] = lfsr[1] ^ lfsr[2] ^ lfsr[4] ^ lfsr[5] ^ lfsr[9] ^ lfsr[11] ^ lfsr[12] ^ lfsr[13] ^ lfsr[18] ^ lfsr[23] ^ lfsr[24] ^ lfsr[29] ^ data_i[1] ^ data_i[2] ^ data_i[4] ^ data_i[5] ^ data_i[9] ^ data_i[11] ^ data_i[12] ^ data_i[13] ^ data_i[18] ^ data_i[23] ^ data_i[24] ^ data_i[29];
   assign lfsr_next[10] = lfsr[0] ^ lfsr[2] ^ lfsr[3] ^ lfsr[5] ^ lfsr[9] ^ lfsr[13] ^ lfsr[14] ^ lfsr[16] ^ lfsr[19] ^ lfsr[26] ^ lfsr[28] ^ lfsr[29] ^ lfsr[31] ^ data_i[0] ^ data_i[2] ^ data_i[3] ^ data_i[5] ^ data_i[9] ^ data_i[13] ^ data_i[14] ^ data_i[16] ^ data_i[19] ^ data_i[26] ^ data_i[28] ^ data_i[29] ^ data_i[31];
   assign lfsr_next[11] = lfsr[0] ^ lfsr[1] ^ lfsr[3] ^ lfsr[4] ^ lfsr[9] ^ lfsr[12] ^ lfsr[14] ^ lfsr[15] ^ lfsr[16] ^ lfsr[17] ^ lfsr[20] ^ lfsr[24] ^ lfsr[25] ^ lfsr[26] ^ lfsr[27] ^ lfsr[28] ^ lfsr[31] ^ data_i[0] ^ data_i[1] ^ data_i[3] ^ data_i[4] ^ data_i[9] ^ data_i[12] ^ data_i[14] ^ data_i[15] ^ data_i[16] ^ data_i[17] ^ data_i[20] ^ data_i[24] ^ data_i[25] ^ data_i[26] ^ data_i[27] ^ data_i[28] ^ data_i[31];
   assign lfsr_next[12] = lfsr[0] ^ lfsr[1] ^ lfsr[2] ^ lfsr[4] ^ lfsr[5] ^ lfsr[6] ^ lfsr[9] ^ lfsr[12] ^ lfsr[13] ^ lfsr[15] ^ lfsr[17] ^ lfsr[18] ^ lfsr[21] ^ lfsr[24] ^ lfsr[27] ^ lfsr[30] ^ lfsr[31] ^ data_i[0] ^ data_i[1] ^ data_i[2] ^ data_i[4] ^ data_i[5] ^ data_i[6] ^ data_i[9] ^ data_i[12] ^ data_i[13] ^ data_i[15] ^ data_i[17] ^ data_i[18] ^ data_i[21] ^ data_i[24] ^ data_i[27] ^ data_i[30] ^ data_i[31];
   assign lfsr_next[13] = lfsr[1] ^ lfsr[2] ^ lfsr[3] ^ lfsr[5] ^ lfsr[6] ^ lfsr[7] ^ lfsr[10] ^ lfsr[13] ^ lfsr[14] ^ lfsr[16] ^ lfsr[18] ^ lfsr[19] ^ lfsr[22] ^ lfsr[25] ^ lfsr[28] ^ lfsr[31] ^ data_i[1] ^ data_i[2] ^ data_i[3] ^ data_i[5] ^ data_i[6] ^ data_i[7] ^ data_i[10] ^ data_i[13] ^ data_i[14] ^ data_i[16] ^ data_i[18] ^ data_i[19] ^ data_i[22] ^ data_i[25] ^ data_i[28] ^ data_i[31];
   assign lfsr_next[14] = lfsr[2] ^ lfsr[3] ^ lfsr[4] ^ lfsr[6] ^ lfsr[7] ^ lfsr[8] ^ lfsr[11] ^ lfsr[14] ^ lfsr[15] ^ lfsr[17] ^ lfsr[19] ^ lfsr[20] ^ lfsr[23] ^ lfsr[26] ^ lfsr[29] ^ data_i[2] ^ data_i[3] ^ data_i[4] ^ data_i[6] ^ data_i[7] ^ data_i[8] ^ data_i[11] ^ data_i[14] ^ data_i[15] ^ data_i[17] ^ data_i[19] ^ data_i[20] ^ data_i[23] ^ data_i[26] ^ data_i[29];
   assign lfsr_next[15] = lfsr[3] ^ lfsr[4] ^ lfsr[5] ^ lfsr[7] ^ lfsr[8] ^ lfsr[9] ^ lfsr[12] ^ lfsr[15] ^ lfsr[16] ^ lfsr[18] ^ lfsr[20] ^ lfsr[21] ^ lfsr[24] ^ lfsr[27] ^ lfsr[30] ^ data_i[3] ^ data_i[4] ^ data_i[5] ^ data_i[7] ^ data_i[8] ^ data_i[9] ^ data_i[12] ^ data_i[15] ^ data_i[16] ^ data_i[18] ^ data_i[20] ^ data_i[21] ^ data_i[24] ^ data_i[27] ^ data_i[30];
   assign lfsr_next[16] = lfsr[0] ^ lfsr[4] ^ lfsr[5] ^ lfsr[8] ^ lfsr[12] ^ lfsr[13] ^ lfsr[17] ^ lfsr[19] ^ lfsr[21] ^ lfsr[22] ^ lfsr[24] ^ lfsr[26] ^ lfsr[29] ^ lfsr[30] ^ data_i[0] ^ data_i[4] ^ data_i[5] ^ data_i[8] ^ data_i[12] ^ data_i[13] ^ data_i[17] ^ data_i[19] ^ data_i[21] ^ data_i[22] ^ data_i[24] ^ data_i[26] ^ data_i[29] ^ data_i[30];
   assign lfsr_next[17] = lfsr[1] ^ lfsr[5] ^ lfsr[6] ^ lfsr[9] ^ lfsr[13] ^ lfsr[14] ^ lfsr[18] ^ lfsr[20] ^ lfsr[22] ^ lfsr[23] ^ lfsr[25] ^ lfsr[27] ^ lfsr[30] ^ lfsr[31] ^ data_i[1] ^ data_i[5] ^ data_i[6] ^ data_i[9] ^ data_i[13] ^ data_i[14] ^ data_i[18] ^ data_i[20] ^ data_i[22] ^ data_i[23] ^ data_i[25] ^ data_i[27] ^ data_i[30] ^ data_i[31];
   assign lfsr_next[18] = lfsr[2] ^ lfsr[6] ^ lfsr[7] ^ lfsr[10] ^ lfsr[14] ^ lfsr[15] ^ lfsr[19] ^ lfsr[21] ^ lfsr[23] ^ lfsr[24] ^ lfsr[26] ^ lfsr[28] ^ lfsr[31] ^ data_i[2] ^ data_i[6] ^ data_i[7] ^ data_i[10] ^ data_i[14] ^ data_i[15] ^ data_i[19] ^ data_i[21] ^ data_i[23] ^ data_i[24] ^ data_i[26] ^ data_i[28] ^ data_i[31];
   assign lfsr_next[19] = lfsr[3] ^ lfsr[7] ^ lfsr[8] ^ lfsr[11] ^ lfsr[15] ^ lfsr[16] ^ lfsr[20] ^ lfsr[22] ^ lfsr[24] ^ lfsr[25] ^ lfsr[27] ^ lfsr[29] ^ data_i[3] ^ data_i[7] ^ data_i[8] ^ data_i[11] ^ data_i[15] ^ data_i[16] ^ data_i[20] ^ data_i[22] ^ data_i[24] ^ data_i[25] ^ data_i[27] ^ data_i[29];
   assign lfsr_next[20] = lfsr[4] ^ lfsr[8] ^ lfsr[9] ^ lfsr[12] ^ lfsr[16] ^ lfsr[17] ^ lfsr[21] ^ lfsr[23] ^ lfsr[25] ^ lfsr[26] ^ lfsr[28] ^ lfsr[30] ^ data_i[4] ^ data_i[8] ^ data_i[9] ^ data_i[12] ^ data_i[16] ^ data_i[17] ^ data_i[21] ^ data_i[23] ^ data_i[25] ^ data_i[26] ^ data_i[28] ^ data_i[30];
   assign lfsr_next[21] = lfsr[5] ^ lfsr[9] ^ lfsr[10] ^ lfsr[13] ^ lfsr[17] ^ lfsr[18] ^ lfsr[22] ^ lfsr[24] ^ lfsr[26] ^ lfsr[27] ^ lfsr[29] ^ lfsr[31] ^ data_i[5] ^ data_i[9] ^ data_i[10] ^ data_i[13] ^ data_i[17] ^ data_i[18] ^ data_i[22] ^ data_i[24] ^ data_i[26] ^ data_i[27] ^ data_i[29] ^ data_i[31];
   assign lfsr_next[22] = lfsr[0] ^ lfsr[9] ^ lfsr[11] ^ lfsr[12] ^ lfsr[14] ^ lfsr[16] ^ lfsr[18] ^ lfsr[19] ^ lfsr[23] ^ lfsr[24] ^ lfsr[26] ^ lfsr[27] ^ lfsr[29] ^ lfsr[31] ^ data_i[0] ^ data_i[9] ^ data_i[11] ^ data_i[12] ^ data_i[14] ^ data_i[16] ^ data_i[18] ^ data_i[19] ^ data_i[23] ^ data_i[24] ^ data_i[26] ^ data_i[27] ^ data_i[29] ^ data_i[31];
   assign lfsr_next[23] = lfsr[0] ^ lfsr[1] ^ lfsr[6] ^ lfsr[9] ^ lfsr[13] ^ lfsr[15] ^ lfsr[16] ^ lfsr[17] ^ lfsr[19] ^ lfsr[20] ^ lfsr[26] ^ lfsr[27] ^ lfsr[29] ^ lfsr[31] ^ data_i[0] ^ data_i[1] ^ data_i[6] ^ data_i[9] ^ data_i[13] ^ data_i[15] ^ data_i[16] ^ data_i[17] ^ data_i[19] ^ data_i[20] ^ data_i[26] ^ data_i[27] ^ data_i[29] ^ data_i[31];
   assign lfsr_next[24] = lfsr[1] ^ lfsr[2] ^ lfsr[7] ^ lfsr[10] ^ lfsr[14] ^ lfsr[16] ^ lfsr[17] ^ lfsr[18] ^ lfsr[20] ^ lfsr[21] ^ lfsr[27] ^ lfsr[28] ^ lfsr[30] ^ data_i[1] ^ data_i[2] ^ data_i[7] ^ data_i[10] ^ data_i[14] ^ data_i[16] ^ data_i[17] ^ data_i[18] ^ data_i[20] ^ data_i[21] ^ data_i[27] ^ data_i[28] ^ data_i[30];
   assign lfsr_next[25] = lfsr[2] ^ lfsr[3] ^ lfsr[8] ^ lfsr[11] ^ lfsr[15] ^ lfsr[17] ^ lfsr[18] ^ lfsr[19] ^ lfsr[21] ^ lfsr[22] ^ lfsr[28] ^ lfsr[29] ^ lfsr[31] ^ data_i[2] ^ data_i[3] ^ data_i[8] ^ data_i[11] ^ data_i[15] ^ data_i[17] ^ data_i[18] ^ data_i[19] ^ data_i[21] ^ data_i[22] ^ data_i[28] ^ data_i[29] ^ data_i[31];
   assign lfsr_next[26] = lfsr[0] ^ lfsr[3] ^ lfsr[4] ^ lfsr[6] ^ lfsr[10] ^ lfsr[18] ^ lfsr[19] ^ lfsr[20] ^ lfsr[22] ^ lfsr[23] ^ lfsr[24] ^ lfsr[25] ^ lfsr[26] ^ lfsr[28] ^ lfsr[31] ^ data_i[0] ^ data_i[3] ^ data_i[4] ^ data_i[6] ^ data_i[10] ^ data_i[18] ^ data_i[19] ^ data_i[20] ^ data_i[22] ^ data_i[23] ^ data_i[24] ^ data_i[25] ^ data_i[26] ^ data_i[28] ^ data_i[31];
   assign lfsr_next[27] = lfsr[1] ^ lfsr[4] ^ lfsr[5] ^ lfsr[7] ^ lfsr[11] ^ lfsr[19] ^ lfsr[20] ^ lfsr[21] ^ lfsr[23] ^ lfsr[24] ^ lfsr[25] ^ lfsr[26] ^ lfsr[27] ^ lfsr[29] ^ data_i[1] ^ data_i[4] ^ data_i[5] ^ data_i[7] ^ data_i[11] ^ data_i[19] ^ data_i[20] ^ data_i[21] ^ data_i[23] ^ data_i[24] ^ data_i[25] ^ data_i[26] ^ data_i[27] ^ data_i[29];
   assign lfsr_next[28] = lfsr[2] ^ lfsr[5] ^ lfsr[6] ^ lfsr[8] ^ lfsr[12] ^ lfsr[20] ^ lfsr[21] ^ lfsr[22] ^ lfsr[24] ^ lfsr[25] ^ lfsr[26] ^ lfsr[27] ^ lfsr[28] ^ lfsr[30] ^ data_i[2] ^ data_i[5] ^ data_i[6] ^ data_i[8] ^ data_i[12] ^ data_i[20] ^ data_i[21] ^ data_i[22] ^ data_i[24] ^ data_i[25] ^ data_i[26] ^ data_i[27] ^ data_i[28] ^ data_i[30];
   assign lfsr_next[29] = lfsr[3] ^ lfsr[6] ^ lfsr[7] ^ lfsr[9] ^ lfsr[13] ^ lfsr[21] ^ lfsr[22] ^ lfsr[23] ^ lfsr[25] ^ lfsr[26] ^ lfsr[27] ^ lfsr[28] ^ lfsr[29] ^ lfsr[31] ^ data_i[3] ^ data_i[6] ^ data_i[7] ^ data_i[9] ^ data_i[13] ^ data_i[21] ^ data_i[22] ^ data_i[23] ^ data_i[25] ^ data_i[26] ^ data_i[27] ^ data_i[28] ^ data_i[29] ^ data_i[31];
   assign lfsr_next[30] = lfsr[4] ^ lfsr[7] ^ lfsr[8] ^ lfsr[10] ^ lfsr[14] ^ lfsr[22] ^ lfsr[23] ^ lfsr[24] ^ lfsr[26] ^ lfsr[27] ^ lfsr[28] ^ lfsr[29] ^ lfsr[30] ^ data_i[4] ^ data_i[7] ^ data_i[8] ^ data_i[10] ^ data_i[14] ^ data_i[22] ^ data_i[23] ^ data_i[24] ^ data_i[26] ^ data_i[27] ^ data_i[28] ^ data_i[29] ^ data_i[30];
   assign lfsr_next[31] = lfsr[5] ^ lfsr[8] ^ lfsr[9] ^ lfsr[11] ^ lfsr[15] ^ lfsr[23] ^ lfsr[24] ^ lfsr[25] ^ lfsr[27] ^ lfsr[28] ^ lfsr[29] ^ lfsr[30] ^ lfsr[31] ^ data_i[5] ^ data_i[8] ^ data_i[9] ^ data_i[11] ^ data_i[15] ^ data_i[23] ^ data_i[24] ^ data_i[25] ^ data_i[27] ^ data_i[28] ^ data_i[29] ^ data_i[30] ^ data_i[31];
 end else if ( DATA_W == 64 ) begin
	assign lfsr_next[0] = lfsr[0] ^ lfsr[2] ^ lfsr[5] ^ lfsr[12] ^ lfsr[13] ^ lfsr[15] ^ lfsr[16] ^ lfsr[18] ^ lfsr[21] ^ lfsr[22] ^ lfsr[23] ^ lfsr[26] ^ lfsr[28] ^ lfsr[29] ^ lfsr[31] ^ data_i[0] ^ data_i[6] ^ data_i[9] ^ data_i[10] ^ data_i[12] ^ data_i[16] ^ data_i[24] ^ data_i[25] ^ data_i[26] ^ data_i[28] ^ data_i[29] ^ data_i[30] ^ data_i[31] ^ data_i[32] ^ data_i[34] ^ data_i[37] ^ data_i[44] ^ data_i[45] ^ data_i[47] ^ data_i[48] ^ data_i[50] ^ data_i[53] ^ data_i[54] ^ data_i[55] ^ data_i[58] ^ data_i[60] ^ data_i[61] ^ data_i[63];
    assign lfsr_next[1] = lfsr[1] ^ lfsr[2] ^ lfsr[3] ^ lfsr[5] ^ lfsr[6] ^ lfsr[12] ^ lfsr[14] ^ lfsr[15] ^ lfsr[17] ^ lfsr[18] ^ lfsr[19] ^ lfsr[21] ^ lfsr[24] ^ lfsr[26] ^ lfsr[27] ^ lfsr[28] ^ lfsr[30] ^ lfsr[31] ^ data_i[0] ^ data_i[1] ^ data_i[6] ^ data_i[7] ^ data_i[9] ^ data_i[11] ^ data_i[12] ^ data_i[13] ^ data_i[16] ^ data_i[17] ^ data_i[24] ^ data_i[27] ^ data_i[28] ^ data_i[33] ^ data_i[34] ^ data_i[35] ^ data_i[37] ^ data_i[38] ^ data_i[44] ^ data_i[46] ^ data_i[47] ^ data_i[49] ^ data_i[50] ^ data_i[51] ^ data_i[53] ^ data_i[56] ^ data_i[58] ^ data_i[59] ^ data_i[60] ^ data_i[62] ^ data_i[63];
    assign lfsr_next[2] = lfsr[0] ^ lfsr[3] ^ lfsr[4] ^ lfsr[5] ^ lfsr[6] ^ lfsr[7] ^ lfsr[12] ^ lfsr[19] ^ lfsr[20] ^ lfsr[21] ^ lfsr[23] ^ lfsr[25] ^ lfsr[26] ^ lfsr[27] ^ data_i[0] ^ data_i[1] ^ data_i[2] ^ data_i[6] ^ data_i[7] ^ data_i[8] ^ data_i[9] ^ data_i[13] ^ data_i[14] ^ data_i[16] ^ data_i[17] ^ data_i[18] ^ data_i[24] ^ data_i[26] ^ data_i[30] ^ data_i[31] ^ data_i[32] ^ data_i[35] ^ data_i[36] ^ data_i[37] ^ data_i[38] ^ data_i[39] ^ data_i[44] ^ data_i[51] ^ data_i[52] ^ data_i[53] ^ data_i[55] ^ data_i[57] ^ data_i[58] ^ data_i[59];
    assign lfsr_next[3] = lfsr[0] ^ lfsr[1] ^ lfsr[4] ^ lfsr[5] ^ lfsr[6] ^ lfsr[7] ^ lfsr[8] ^ lfsr[13] ^ lfsr[20] ^ lfsr[21] ^ lfsr[22] ^ lfsr[24] ^ lfsr[26] ^ lfsr[27] ^ lfsr[28] ^ data_i[1] ^ data_i[2] ^ data_i[3] ^ data_i[7] ^ data_i[8] ^ data_i[9] ^ data_i[10] ^ data_i[14] ^ data_i[15] ^ data_i[17] ^ data_i[18] ^ data_i[19] ^ data_i[25] ^ data_i[27] ^ data_i[31] ^ data_i[32] ^ data_i[33] ^ data_i[36] ^ data_i[37] ^ data_i[38] ^ data_i[39] ^ data_i[40] ^ data_i[45] ^ data_i[52] ^ data_i[53] ^ data_i[54] ^ data_i[56] ^ data_i[58] ^ data_i[59] ^ data_i[60];
    assign lfsr_next[4] = lfsr[1] ^ lfsr[6] ^ lfsr[7] ^ lfsr[8] ^ lfsr[9] ^ lfsr[12] ^ lfsr[13] ^ lfsr[14] ^ lfsr[15] ^ lfsr[16] ^ lfsr[18] ^ lfsr[25] ^ lfsr[26] ^ lfsr[27] ^ lfsr[31] ^ data_i[0] ^ data_i[2] ^ data_i[3] ^ data_i[4] ^ data_i[6] ^ data_i[8] ^ data_i[11] ^ data_i[12] ^ data_i[15] ^ data_i[18] ^ data_i[19] ^ data_i[20] ^ data_i[24] ^ data_i[25] ^ data_i[29] ^ data_i[30] ^ data_i[31] ^ data_i[33] ^ data_i[38] ^ data_i[39] ^ data_i[40] ^ data_i[41] ^ data_i[44] ^ data_i[45] ^ data_i[46] ^ data_i[47] ^ data_i[48] ^ data_i[50] ^ data_i[57] ^ data_i[58] ^ data_i[59] ^ data_i[63];
    assign lfsr_next[5] = lfsr[5] ^ lfsr[7] ^ lfsr[8] ^ lfsr[9] ^ lfsr[10] ^ lfsr[12] ^ lfsr[14] ^ lfsr[17] ^ lfsr[18] ^ lfsr[19] ^ lfsr[21] ^ lfsr[22] ^ lfsr[23] ^ lfsr[27] ^ lfsr[29] ^ lfsr[31] ^ data_i[0] ^ data_i[1] ^ data_i[3] ^ data_i[4] ^ data_i[5] ^ data_i[6] ^ data_i[7] ^ data_i[10] ^ data_i[13] ^ data_i[19] ^ data_i[20] ^ data_i[21] ^ data_i[24] ^ data_i[28] ^ data_i[29] ^ data_i[37] ^ data_i[39] ^ data_i[40] ^ data_i[41] ^ data_i[42] ^ data_i[44] ^ data_i[46] ^ data_i[49] ^ data_i[50] ^ data_i[51] ^ data_i[53] ^ data_i[54] ^ data_i[55] ^ data_i[59] ^ data_i[61] ^ data_i[63];
    assign lfsr_next[6] = lfsr[6] ^ lfsr[8] ^ lfsr[9] ^ lfsr[10] ^ lfsr[11] ^ lfsr[13] ^ lfsr[15] ^ lfsr[18] ^ lfsr[19] ^ lfsr[20] ^ lfsr[22] ^ lfsr[23] ^ lfsr[24] ^ lfsr[28] ^ lfsr[30] ^ data_i[1] ^ data_i[2] ^ data_i[4] ^ data_i[5] ^ data_i[6] ^ data_i[7] ^ data_i[8] ^ data_i[11] ^ data_i[14] ^ data_i[20] ^ data_i[21] ^ data_i[22] ^ data_i[25] ^ data_i[29] ^ data_i[30] ^ data_i[38] ^ data_i[40] ^ data_i[41] ^ data_i[42] ^ data_i[43] ^ data_i[45] ^ data_i[47] ^ data_i[50] ^ data_i[51] ^ data_i[52] ^ data_i[54] ^ data_i[55] ^ data_i[56] ^ data_i[60] ^ data_i[62];
    assign lfsr_next[7] = lfsr[0] ^ lfsr[2] ^ lfsr[5] ^ lfsr[7] ^ lfsr[9] ^ lfsr[10] ^ lfsr[11] ^ lfsr[13] ^ lfsr[14] ^ lfsr[15] ^ lfsr[18] ^ lfsr[19] ^ lfsr[20] ^ lfsr[22] ^ lfsr[24] ^ lfsr[25] ^ lfsr[26] ^ lfsr[28] ^ data_i[0] ^ data_i[2] ^ data_i[3] ^ data_i[5] ^ data_i[7] ^ data_i[8] ^ data_i[10] ^ data_i[15] ^ data_i[16] ^ data_i[21] ^ data_i[22] ^ data_i[23] ^ data_i[24] ^ data_i[25] ^ data_i[28] ^ data_i[29] ^ data_i[32] ^ data_i[34] ^ data_i[37] ^ data_i[39] ^ data_i[41] ^ data_i[42] ^ data_i[43] ^ data_i[45] ^ data_i[46] ^ data_i[47] ^ data_i[50] ^ data_i[51] ^ data_i[52] ^ data_i[54] ^ data_i[56] ^ data_i[57] ^ data_i[58] ^ data_i[60];
    assign lfsr_next[8] = lfsr[0] ^ lfsr[1] ^ lfsr[2] ^ lfsr[3] ^ lfsr[5] ^ lfsr[6] ^ lfsr[8] ^ lfsr[10] ^ lfsr[11] ^ lfsr[13] ^ lfsr[14] ^ lfsr[18] ^ lfsr[19] ^ lfsr[20] ^ lfsr[22] ^ lfsr[25] ^ lfsr[27] ^ lfsr[28] ^ lfsr[31] ^ data_i[0] ^ data_i[1] ^ data_i[3] ^ data_i[4] ^ data_i[8] ^ data_i[10] ^ data_i[11] ^ data_i[12] ^ data_i[17] ^ data_i[22] ^ data_i[23] ^ data_i[28] ^ data_i[31] ^ data_i[32] ^ data_i[33] ^ data_i[34] ^ data_i[35] ^ data_i[37] ^ data_i[38] ^ data_i[40] ^ data_i[42] ^ data_i[43] ^ data_i[45] ^ data_i[46] ^ data_i[50] ^ data_i[51] ^ data_i[52] ^ data_i[54] ^ data_i[57] ^ data_i[59] ^ data_i[60] ^ data_i[63];
    assign lfsr_next[9] = lfsr[0] ^ lfsr[1] ^ lfsr[2] ^ lfsr[3] ^ lfsr[4] ^ lfsr[6] ^ lfsr[7] ^ lfsr[9] ^ lfsr[11] ^ lfsr[12] ^ lfsr[14] ^ lfsr[15] ^ lfsr[19] ^ lfsr[20] ^ lfsr[21] ^ lfsr[23] ^ lfsr[26] ^ lfsr[28] ^ lfsr[29] ^ data_i[1] ^ data_i[2] ^ data_i[4] ^ data_i[5] ^ data_i[9] ^ data_i[11] ^ data_i[12] ^ data_i[13] ^ data_i[18] ^ data_i[23] ^ data_i[24] ^ data_i[29] ^ data_i[32] ^ data_i[33] ^ data_i[34] ^ data_i[35] ^ data_i[36] ^ data_i[38] ^ data_i[39] ^ data_i[41] ^ data_i[43] ^ data_i[44] ^ data_i[46] ^ data_i[47] ^ data_i[51] ^ data_i[52] ^ data_i[53] ^ data_i[55] ^ data_i[58] ^ data_i[60] ^ data_i[61];
    assign lfsr_next[10] = lfsr[0] ^ lfsr[1] ^ lfsr[3] ^ lfsr[4] ^ lfsr[7] ^ lfsr[8] ^ lfsr[10] ^ lfsr[18] ^ lfsr[20] ^ lfsr[23] ^ lfsr[24] ^ lfsr[26] ^ lfsr[27] ^ lfsr[28] ^ lfsr[30] ^ lfsr[31] ^ data_i[0] ^ data_i[2] ^ data_i[3] ^ data_i[5] ^ data_i[9] ^ data_i[13] ^ data_i[14] ^ data_i[16] ^ data_i[19] ^ data_i[26] ^ data_i[28] ^ data_i[29] ^ data_i[31] ^ data_i[32] ^ data_i[33] ^ data_i[35] ^ data_i[36] ^ data_i[39] ^ data_i[40] ^ data_i[42] ^ data_i[50] ^ data_i[52] ^ data_i[55] ^ data_i[56] ^ data_i[58] ^ data_i[59] ^ data_i[60] ^ data_i[62] ^ data_i[63];
    assign lfsr_next[11] = lfsr[1] ^ lfsr[4] ^ lfsr[8] ^ lfsr[9] ^ lfsr[11] ^ lfsr[12] ^ lfsr[13] ^ lfsr[15] ^ lfsr[16] ^ lfsr[18] ^ lfsr[19] ^ lfsr[22] ^ lfsr[23] ^ lfsr[24] ^ lfsr[25] ^ lfsr[26] ^ lfsr[27] ^ data_i[0] ^ data_i[1] ^ data_i[3] ^ data_i[4] ^ data_i[9] ^ data_i[12] ^ data_i[14] ^ data_i[15] ^ data_i[16] ^ data_i[17] ^ data_i[20] ^ data_i[24] ^ data_i[25] ^ data_i[26] ^ data_i[27] ^ data_i[28] ^ data_i[31] ^ data_i[33] ^ data_i[36] ^ data_i[40] ^ data_i[41] ^ data_i[43] ^ data_i[44] ^ data_i[45] ^ data_i[47] ^ data_i[48] ^ data_i[50] ^ data_i[51] ^ data_i[54] ^ data_i[55] ^ data_i[56] ^ data_i[57] ^ data_i[58] ^ data_i[59];
    assign lfsr_next[12] = lfsr[9] ^ lfsr[10] ^ lfsr[14] ^ lfsr[15] ^ lfsr[17] ^ lfsr[18] ^ lfsr[19] ^ lfsr[20] ^ lfsr[21] ^ lfsr[22] ^ lfsr[24] ^ lfsr[25] ^ lfsr[27] ^ lfsr[29] ^ lfsr[31] ^ data_i[0] ^ data_i[1] ^ data_i[2] ^ data_i[4] ^ data_i[5] ^ data_i[6] ^ data_i[9] ^ data_i[12] ^ data_i[13] ^ data_i[15] ^ data_i[17] ^ data_i[18] ^ data_i[21] ^ data_i[24] ^ data_i[27] ^ data_i[30] ^ data_i[31] ^ data_i[41] ^ data_i[42] ^ data_i[46] ^ data_i[47] ^ data_i[49] ^ data_i[50] ^ data_i[51] ^ data_i[52] ^ data_i[53] ^ data_i[54] ^ data_i[56] ^ data_i[57] ^ data_i[59] ^ data_i[61] ^ data_i[63];
    assign lfsr_next[13] = lfsr[0] ^ lfsr[10] ^ lfsr[11] ^ lfsr[15] ^ lfsr[16] ^ lfsr[18] ^ lfsr[19] ^ lfsr[20] ^ lfsr[21] ^ lfsr[22] ^ lfsr[23] ^ lfsr[25] ^ lfsr[26] ^ lfsr[28] ^ lfsr[30] ^ data_i[1] ^ data_i[2] ^ data_i[3] ^ data_i[5] ^ data_i[6] ^ data_i[7] ^ data_i[10] ^ data_i[13] ^ data_i[14] ^ data_i[16] ^ data_i[18] ^ data_i[19] ^ data_i[22] ^ data_i[25] ^ data_i[28] ^ data_i[31] ^ data_i[32] ^ data_i[42] ^ data_i[43] ^ data_i[47] ^ data_i[48] ^ data_i[50] ^ data_i[51] ^ data_i[52] ^ data_i[53] ^ data_i[54] ^ data_i[55] ^ data_i[57] ^ data_i[58] ^ data_i[60] ^ data_i[62];
    assign lfsr_next[14] = lfsr[0] ^ lfsr[1] ^ lfsr[11] ^ lfsr[12] ^ lfsr[16] ^ lfsr[17] ^ lfsr[19] ^ lfsr[20] ^ lfsr[21] ^ lfsr[22] ^ lfsr[23] ^ lfsr[24] ^ lfsr[26] ^ lfsr[27] ^ lfsr[29] ^ lfsr[31] ^ data_i[2] ^ data_i[3] ^ data_i[4] ^ data_i[6] ^ data_i[7] ^ data_i[8] ^ data_i[11] ^ data_i[14] ^ data_i[15] ^ data_i[17] ^ data_i[19] ^ data_i[20] ^ data_i[23] ^ data_i[26] ^ data_i[29] ^ data_i[32] ^ data_i[33] ^ data_i[43] ^ data_i[44] ^ data_i[48] ^ data_i[49] ^ data_i[51] ^ data_i[52] ^ data_i[53] ^ data_i[54] ^ data_i[55] ^ data_i[56] ^ data_i[58] ^ data_i[59] ^ data_i[61] ^ data_i[63];
    assign lfsr_next[15] = lfsr[1] ^ lfsr[2] ^ lfsr[12] ^ lfsr[13] ^ lfsr[17] ^ lfsr[18] ^ lfsr[20] ^ lfsr[21] ^ lfsr[22] ^ lfsr[23] ^ lfsr[24] ^ lfsr[25] ^ lfsr[27] ^ lfsr[28] ^ lfsr[30] ^ data_i[3] ^ data_i[4] ^ data_i[5] ^ data_i[7] ^ data_i[8] ^ data_i[9] ^ data_i[12] ^ data_i[15] ^ data_i[16] ^ data_i[18] ^ data_i[20] ^ data_i[21] ^ data_i[24] ^ data_i[27] ^ data_i[30] ^ data_i[33] ^ data_i[34] ^ data_i[44] ^ data_i[45] ^ data_i[49] ^ data_i[50] ^ data_i[52] ^ data_i[53] ^ data_i[54] ^ data_i[55] ^ data_i[56] ^ data_i[57] ^ data_i[59] ^ data_i[60] ^ data_i[62];
    assign lfsr_next[16] = lfsr[0] ^ lfsr[3] ^ lfsr[5] ^ lfsr[12] ^ lfsr[14] ^ lfsr[15] ^ lfsr[16] ^ lfsr[19] ^ lfsr[24] ^ lfsr[25] ^ data_i[0] ^ data_i[4] ^ data_i[5] ^ data_i[8] ^ data_i[12] ^ data_i[13] ^ data_i[17] ^ data_i[19] ^ data_i[21] ^ data_i[22] ^ data_i[24] ^ data_i[26] ^ data_i[29] ^ data_i[30] ^ data_i[32] ^ data_i[35] ^ data_i[37] ^ data_i[44] ^ data_i[46] ^ data_i[47] ^ data_i[48] ^ data_i[51] ^ data_i[56] ^ data_i[57];
    assign lfsr_next[17] = lfsr[1] ^ lfsr[4] ^ lfsr[6] ^ lfsr[13] ^ lfsr[15] ^ lfsr[16] ^ lfsr[17] ^ lfsr[20] ^ lfsr[25] ^ lfsr[26] ^ data_i[1] ^ data_i[5] ^ data_i[6] ^ data_i[9] ^ data_i[13] ^ data_i[14] ^ data_i[18] ^ data_i[20] ^ data_i[22] ^ data_i[23] ^ data_i[25] ^ data_i[27] ^ data_i[30] ^ data_i[31] ^ data_i[33] ^ data_i[36] ^ data_i[38] ^ data_i[45] ^ data_i[47] ^ data_i[48] ^ data_i[49] ^ data_i[52] ^ data_i[57] ^ data_i[58];
    assign lfsr_next[18] = lfsr[0] ^ lfsr[2] ^ lfsr[5] ^ lfsr[7] ^ lfsr[14] ^ lfsr[16] ^ lfsr[17] ^ lfsr[18] ^ lfsr[21] ^ lfsr[26] ^ lfsr[27] ^ data_i[2] ^ data_i[6] ^ data_i[7] ^ data_i[10] ^ data_i[14] ^ data_i[15] ^ data_i[19] ^ data_i[21] ^ data_i[23] ^ data_i[24] ^ data_i[26] ^ data_i[28] ^ data_i[31] ^ data_i[32] ^ data_i[34] ^ data_i[37] ^ data_i[39] ^ data_i[46] ^ data_i[48] ^ data_i[49] ^ data_i[50] ^ data_i[53] ^ data_i[58] ^ data_i[59];
    assign lfsr_next[19] = lfsr[0] ^ lfsr[1] ^ lfsr[3] ^ lfsr[6] ^ lfsr[8] ^ lfsr[15] ^ lfsr[17] ^ lfsr[18] ^ lfsr[19] ^ lfsr[22] ^ lfsr[27] ^ lfsr[28] ^ data_i[3] ^ data_i[7] ^ data_i[8] ^ data_i[11] ^ data_i[15] ^ data_i[16] ^ data_i[20] ^ data_i[22] ^ data_i[24] ^ data_i[25] ^ data_i[27] ^ data_i[29] ^ data_i[32] ^ data_i[33] ^ data_i[35] ^ data_i[38] ^ data_i[40] ^ data_i[47] ^ data_i[49] ^ data_i[50] ^ data_i[51] ^ data_i[54] ^ data_i[59] ^ data_i[60];
    assign lfsr_next[20] = lfsr[1] ^ lfsr[2] ^ lfsr[4] ^ lfsr[7] ^ lfsr[9] ^ lfsr[16] ^ lfsr[18] ^ lfsr[19] ^ lfsr[20] ^ lfsr[23] ^ lfsr[28] ^ lfsr[29] ^ data_i[4] ^ data_i[8] ^ data_i[9] ^ data_i[12] ^ data_i[16] ^ data_i[17] ^ data_i[21] ^ data_i[23] ^ data_i[25] ^ data_i[26] ^ data_i[28] ^ data_i[30] ^ data_i[33] ^ data_i[34] ^ data_i[36] ^ data_i[39] ^ data_i[41] ^ data_i[48] ^ data_i[50] ^ data_i[51] ^ data_i[52] ^ data_i[55] ^ data_i[60] ^ data_i[61];
    assign lfsr_next[21] = lfsr[2] ^ lfsr[3] ^ lfsr[5] ^ lfsr[8] ^ lfsr[10] ^ lfsr[17] ^ lfsr[19] ^ lfsr[20] ^ lfsr[21] ^ lfsr[24] ^ lfsr[29] ^ lfsr[30] ^ data_i[5] ^ data_i[9] ^ data_i[10] ^ data_i[13] ^ data_i[17] ^ data_i[18] ^ data_i[22] ^ data_i[24] ^ data_i[26] ^ data_i[27] ^ data_i[29] ^ data_i[31] ^ data_i[34] ^ data_i[35] ^ data_i[37] ^ data_i[40] ^ data_i[42] ^ data_i[49] ^ data_i[51] ^ data_i[52] ^ data_i[53] ^ data_i[56] ^ data_i[61] ^ data_i[62];
    assign lfsr_next[22] = lfsr[2] ^ lfsr[3] ^ lfsr[4] ^ lfsr[5] ^ lfsr[6] ^ lfsr[9] ^ lfsr[11] ^ lfsr[12] ^ lfsr[13] ^ lfsr[15] ^ lfsr[16] ^ lfsr[20] ^ lfsr[23] ^ lfsr[25] ^ lfsr[26] ^ lfsr[28] ^ lfsr[29] ^ lfsr[30] ^ data_i[0] ^ data_i[9] ^ data_i[11] ^ data_i[12] ^ data_i[14] ^ data_i[16] ^ data_i[18] ^ data_i[19] ^ data_i[23] ^ data_i[24] ^ data_i[26] ^ data_i[27] ^ data_i[29] ^ data_i[31] ^ data_i[34] ^ data_i[35] ^ data_i[36] ^ data_i[37] ^ data_i[38] ^ data_i[41] ^ data_i[43] ^ data_i[44] ^ data_i[45] ^ data_i[47] ^ data_i[48] ^ data_i[52] ^ data_i[55] ^ data_i[57] ^ data_i[58] ^ data_i[60] ^ data_i[61] ^ data_i[62];
    assign lfsr_next[23] = lfsr[2] ^ lfsr[3] ^ lfsr[4] ^ lfsr[6] ^ lfsr[7] ^ lfsr[10] ^ lfsr[14] ^ lfsr[15] ^ lfsr[17] ^ lfsr[18] ^ lfsr[22] ^ lfsr[23] ^ lfsr[24] ^ lfsr[27] ^ lfsr[28] ^ lfsr[30] ^ data_i[0] ^ data_i[1] ^ data_i[6] ^ data_i[9] ^ data_i[13] ^ data_i[15] ^ data_i[16] ^ data_i[17] ^ data_i[19] ^ data_i[20] ^ data_i[26] ^ data_i[27] ^ data_i[29] ^ data_i[31] ^ data_i[34] ^ data_i[35] ^ data_i[36] ^ data_i[38] ^ data_i[39] ^ data_i[42] ^ data_i[46] ^ data_i[47] ^ data_i[49] ^ data_i[50] ^ data_i[54] ^ data_i[55] ^ data_i[56] ^ data_i[59] ^ data_i[60] ^ data_i[62];
    assign lfsr_next[24] = lfsr[0] ^ lfsr[3] ^ lfsr[4] ^ lfsr[5] ^ lfsr[7] ^ lfsr[8] ^ lfsr[11] ^ lfsr[15] ^ lfsr[16] ^ lfsr[18] ^ lfsr[19] ^ lfsr[23] ^ lfsr[24] ^ lfsr[25] ^ lfsr[28] ^ lfsr[29] ^ lfsr[31] ^ data_i[1] ^ data_i[2] ^ data_i[7] ^ data_i[10] ^ data_i[14] ^ data_i[16] ^ data_i[17] ^ data_i[18] ^ data_i[20] ^ data_i[21] ^ data_i[27] ^ data_i[28] ^ data_i[30] ^ data_i[32] ^ data_i[35] ^ data_i[36] ^ data_i[37] ^ data_i[39] ^ data_i[40] ^ data_i[43] ^ data_i[47] ^ data_i[48] ^ data_i[50] ^ data_i[51] ^ data_i[55] ^ data_i[56] ^ data_i[57] ^ data_i[60] ^ data_i[61] ^ data_i[63];
    assign lfsr_next[25] = lfsr[1] ^ lfsr[4] ^ lfsr[5] ^ lfsr[6] ^ lfsr[8] ^ lfsr[9] ^ lfsr[12] ^ lfsr[16] ^ lfsr[17] ^ lfsr[19] ^ lfsr[20] ^ lfsr[24] ^ lfsr[25] ^ lfsr[26] ^ lfsr[29] ^ lfsr[30] ^ data_i[2] ^ data_i[3] ^ data_i[8] ^ data_i[11] ^ data_i[15] ^ data_i[17] ^ data_i[18] ^ data_i[19] ^ data_i[21] ^ data_i[22] ^ data_i[28] ^ data_i[29] ^ data_i[31] ^ data_i[33] ^ data_i[36] ^ data_i[37] ^ data_i[38] ^ data_i[40] ^ data_i[41] ^ data_i[44] ^ data_i[48] ^ data_i[49] ^ data_i[51] ^ data_i[52] ^ data_i[56] ^ data_i[57] ^ data_i[58] ^ data_i[61] ^ data_i[62];
    assign lfsr_next[26] = lfsr[6] ^ lfsr[7] ^ lfsr[9] ^ lfsr[10] ^ lfsr[12] ^ lfsr[15] ^ lfsr[16] ^ lfsr[17] ^ lfsr[20] ^ lfsr[22] ^ lfsr[23] ^ lfsr[25] ^ lfsr[27] ^ lfsr[28] ^ lfsr[29] ^ lfsr[30] ^ data_i[0] ^ data_i[3] ^ data_i[4] ^ data_i[6] ^ data_i[10] ^ data_i[18] ^ data_i[19] ^ data_i[20] ^ data_i[22] ^ data_i[23] ^ data_i[24] ^ data_i[25] ^ data_i[26] ^ data_i[28] ^ data_i[31] ^ data_i[38] ^ data_i[39] ^ data_i[41] ^ data_i[42] ^ data_i[44] ^ data_i[47] ^ data_i[48] ^ data_i[49] ^ data_i[52] ^ data_i[54] ^ data_i[55] ^ data_i[57] ^ data_i[59] ^ data_i[60] ^ data_i[61] ^ data_i[62];
    assign lfsr_next[27] = lfsr[0] ^ lfsr[7] ^ lfsr[8] ^ lfsr[10] ^ lfsr[11] ^ lfsr[13] ^ lfsr[16] ^ lfsr[17] ^ lfsr[18] ^ lfsr[21] ^ lfsr[23] ^ lfsr[24] ^ lfsr[26] ^ lfsr[28] ^ lfsr[29] ^ lfsr[30] ^ lfsr[31] ^ data_i[1] ^ data_i[4] ^ data_i[5] ^ data_i[7] ^ data_i[11] ^ data_i[19] ^ data_i[20] ^ data_i[21] ^ data_i[23] ^ data_i[24] ^ data_i[25] ^ data_i[26] ^ data_i[27] ^ data_i[29] ^ data_i[32] ^ data_i[39] ^ data_i[40] ^ data_i[42] ^ data_i[43] ^ data_i[45] ^ data_i[48] ^ data_i[49] ^ data_i[50] ^ data_i[53] ^ data_i[55] ^ data_i[56] ^ data_i[58] ^ data_i[60] ^ data_i[61] ^ data_i[62] ^ data_i[63];
    assign lfsr_next[28] = lfsr[1] ^ lfsr[8] ^ lfsr[9] ^ lfsr[11] ^ lfsr[12] ^ lfsr[14] ^ lfsr[17] ^ lfsr[18] ^ lfsr[19] ^ lfsr[22] ^ lfsr[24] ^ lfsr[25] ^ lfsr[27] ^ lfsr[29] ^ lfsr[30] ^ lfsr[31] ^ data_i[2] ^ data_i[5] ^ data_i[6] ^ data_i[8] ^ data_i[12] ^ data_i[20] ^ data_i[21] ^ data_i[22] ^ data_i[24] ^ data_i[25] ^ data_i[26] ^ data_i[27] ^ data_i[28] ^ data_i[30] ^ data_i[33] ^ data_i[40] ^ data_i[41] ^ data_i[43] ^ data_i[44] ^ data_i[46] ^ data_i[49] ^ data_i[50] ^ data_i[51] ^ data_i[54] ^ data_i[56] ^ data_i[57] ^ data_i[59] ^ data_i[61] ^ data_i[62] ^ data_i[63];
    assign lfsr_next[29] = lfsr[2] ^ lfsr[9] ^ lfsr[10] ^ lfsr[12] ^ lfsr[13] ^ lfsr[15] ^ lfsr[18] ^ lfsr[19] ^ lfsr[20] ^ lfsr[23] ^ lfsr[25] ^ lfsr[26] ^ lfsr[28] ^ lfsr[30] ^ lfsr[31] ^ data_i[3] ^ data_i[6] ^ data_i[7] ^ data_i[9] ^ data_i[13] ^ data_i[21] ^ data_i[22] ^ data_i[23] ^ data_i[25] ^ data_i[26] ^ data_i[27] ^ data_i[28] ^ data_i[29] ^ data_i[31] ^ data_i[34] ^ data_i[41] ^ data_i[42] ^ data_i[44] ^ data_i[45] ^ data_i[47] ^ data_i[50] ^ data_i[51] ^ data_i[52] ^ data_i[55] ^ data_i[57] ^ data_i[58] ^ data_i[60] ^ data_i[62] ^ data_i[63];
    assign lfsr_next[30] = lfsr[0] ^ lfsr[3] ^ lfsr[10] ^ lfsr[11] ^ lfsr[13] ^ lfsr[14] ^ lfsr[16] ^ lfsr[19] ^ lfsr[20] ^ lfsr[21] ^ lfsr[24] ^ lfsr[26] ^ lfsr[27] ^ lfsr[29] ^ lfsr[31] ^ data_i[4] ^ data_i[7] ^ data_i[8] ^ data_i[10] ^ data_i[14] ^ data_i[22] ^ data_i[23] ^ data_i[24] ^ data_i[26] ^ data_i[27] ^ data_i[28] ^ data_i[29] ^ data_i[30] ^ data_i[32] ^ data_i[35] ^ data_i[42] ^ data_i[43] ^ data_i[45] ^ data_i[46] ^ data_i[48] ^ data_i[51] ^ data_i[52] ^ data_i[53] ^ data_i[56] ^ data_i[58] ^ data_i[59] ^ data_i[61] ^ data_i[63];
    assign lfsr_next[31] = lfsr[1] ^ lfsr[4] ^ lfsr[11] ^ lfsr[12] ^ lfsr[14] ^ lfsr[15] ^ lfsr[17] ^ lfsr[20] ^ lfsr[21] ^ lfsr[22] ^ lfsr[25] ^ lfsr[27] ^ lfsr[28] ^ lfsr[30] ^ data_i[5] ^ data_i[8] ^ data_i[9] ^ data_i[11] ^ data_i[15] ^ data_i[23] ^ data_i[24] ^ data_i[25] ^ data_i[27] ^ data_i[28] ^ data_i[29] ^ data_i[30] ^ data_i[31] ^ data_i[33] ^ data_i[36] ^ data_i[43] ^ data_i[44] ^ data_i[46] ^ data_i[47] ^ data_i[49] ^ data_i[52] ^ data_i[53] ^ data_i[54] ^ data_i[57] ^ data_i[59] ^ data_i[60] ^ data_i[62];
end

  always @(posedge clk) begin
    if ( valid_i )  begin
      lfsr_q <= lfsr_next;
    end
  end // always
endmodule // crc
